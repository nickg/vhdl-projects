library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.debugtools.all;

--
entity charrom is
port (Clk : in std_logic;
        address : in integer range 0 to 4095;
        -- chip select, active low       
        cs : in std_logic;
        data_o : out std_logic_vector(7 downto 0);

        writeclk : in std_logic;
        -- Yes, we do have a write enable, because we allow modification of ROMs
        -- in the running machine, unless purposely disabled.  This gives us
        -- something like the WOM that the Amiga had.
        writecs : in std_logic;
        we : in std_logic;
        writeaddress : in unsigned(11 downto 0);
        data_i : in std_logic_vector(7 downto 0)
      );
end charrom;

architecture Behavioral of charrom is

-- 4K x 8bit pre-initialised RAM for character ROM

type ram_t is array (0 to 4095) of std_logic_vector(7 downto 0);
signal ram : ram_t := (

x"3c",x"66",x"6e",x"6e",x"60",x"66",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ ** *** ]
-- [ ** *** ]
-- [ **     ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"3c",x"66",x"66",x"7e",x"66",x"66",x"66",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"7c",x"66",x"66",x"7c",x"66",x"66",x"7e",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"3c",x"66",x"66",x"60",x"60",x"66",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **     ]
-- [ **     ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"7c",x"66",x"66",x"66",x"66",x"66",x"7c",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"7e",x"66",x"60",x"78",x"60",x"66",x"7e",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [ **     ]
-- [ ****   ]
-- [ **     ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"7e",x"66",x"60",x"78",x"60",x"60",x"60",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [ **     ]
-- [ ****   ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [        ]
x"3e",x"66",x"60",x"6e",x"66",x"66",x"3e",x"00",
-- [  ***** ]
-- [ **  ** ]
-- [ **     ]
-- [ ** *** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"66",x"66",x"66",x"7e",x"66",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"7e",x"18",x"18",x"18",x"18",x"18",x"7e",x"00",
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [ ****** ]
-- [        ]
x"7e",x"66",x"06",x"06",x"66",x"66",x"7c",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [     ** ]
-- [     ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"66",x"66",x"6c",x"78",x"6c",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ ** **  ]
-- [ ****   ]
-- [ ** **  ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"60",x"60",x"60",x"60",x"60",x"66",x"7e",x"00",
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"63",x"77",x"7f",x"7f",x"6b",x"63",x"63",x"00",
-- [ **   **]
-- [ *** ***]
-- [ *******]
-- [ *******]
-- [ ** * **]
-- [ **   **]
-- [ **   **]
-- [        ]
x"66",x"66",x"76",x"7e",x"6e",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ *** ** ]
-- [ ****** ]
-- [ ** *** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"3c",x"66",x"66",x"66",x"66",x"66",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"7c",x"66",x"66",x"7e",x"60",x"60",x"60",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [        ]
x"3c",x"66",x"66",x"66",x"6a",x"6c",x"36",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ** * * ]
-- [ ** **  ]
-- [  ** ** ]
-- [        ]
x"7c",x"66",x"66",x"7c",x"66",x"66",x"66",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"3e",x"60",x"70",x"3c",x"0e",x"0e",x"7c",x"00",
-- [  ***** ]
-- [ **     ]
-- [ ***    ]
-- [  ****  ]
-- [    *** ]
-- [    *** ]
-- [ *****  ]
-- [        ]
x"7e",x"18",x"18",x"18",x"18",x"18",x"18",x"00",
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"66",x"66",x"66",x"66",x"66",x"6e",x"3c",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ** *** ]
-- [  ****  ]
-- [        ]
x"66",x"66",x"66",x"2c",x"3c",x"18",x"18",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  * **  ]
-- [  ****  ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"63",x"63",x"6b",x"7f",x"7f",x"77",x"63",x"00",
-- [ **   **]
-- [ **   **]
-- [ ** * **]
-- [ *******]
-- [ *******]
-- [ *** ***]
-- [ **   **]
-- [        ]
x"66",x"66",x"3c",x"18",x"3c",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [  ****  ]
-- [   **   ]
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"66",x"66",x"6e",x"3c",x"18",x"18",x"18",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ ** *** ]
-- [  ****  ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"7e",x"66",x"0c",x"18",x"30",x"76",x"7e",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ *** ** ]
-- [ ****** ]
-- [        ]
x"3c",x"30",x"30",x"30",x"30",x"30",x"3c",x"00",
-- [  ****  ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  ****  ]
-- [        ]
x"3c",x"66",x"60",x"78",x"30",x"30",x"7e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **     ]
-- [ ****   ]
-- [  **    ]
-- [  **    ]
-- [ ****** ]
-- [        ]
x"3c",x"0c",x"0c",x"0c",x"0c",x"0c",x"3c",x"00",
-- [  ****  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [  ****  ]
-- [        ]
x"08",x"1c",x"3e",x"1c",x"1c",x"1c",x"1c",x"00",
-- [    *   ]
-- [   ***  ]
-- [  ***** ]
-- [   ***  ]
-- [   ***  ]
-- [   ***  ]
-- [   ***  ]
-- [        ]
x"00",x"10",x"3f",x"7f",x"3f",x"10",x"00",x"00",
-- [        ]
-- [   *    ]
-- [  ******]
-- [ *******]
-- [  ******]
-- [   *    ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"38",x"38",x"38",x"38",x"38",x"00",x"38",x"00",
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [        ]
-- [  ***   ]
-- [        ]
x"6c",x"6c",x"48",x"00",x"00",x"00",x"00",x"00",
-- [ ** **  ]
-- [ ** **  ]
-- [ *  *   ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"18",x"7e",x"60",x"7e",x"06",x"7e",x"18",x"00",
-- [   **   ]
-- [ ****** ]
-- [ **     ]
-- [ ****** ]
-- [     ** ]
-- [ ****** ]
-- [   **   ]
-- [        ]
x"62",x"66",x"0c",x"18",x"30",x"66",x"46",x"00",
-- [ **   * ]
-- [ **  ** ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ **  ** ]
-- [ *   ** ]
-- [        ]
x"3c",x"66",x"66",x"3c",x"74",x"6e",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ****  ]
-- [ *** *  ]
-- [ ** *** ]
-- [  ***** ]
-- [        ]
x"18",x"18",x"10",x"00",x"00",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   *    ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"1c",x"30",x"30",x"30",x"30",x"30",x"1c",x"00",
-- [   ***  ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [   ***  ]
-- [        ]
x"38",x"0c",x"0c",x"0c",x"0c",x"0c",x"38",x"00",
-- [  ***   ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [  ***   ]
-- [        ]
x"08",x"2a",x"1c",x"7f",x"1c",x"2a",x"08",x"00",
-- [    *   ]
-- [  * * * ]
-- [   ***  ]
-- [ *******]
-- [   ***  ]
-- [  * * * ]
-- [    *   ]
-- [        ]
x"00",x"18",x"18",x"7e",x"18",x"18",x"00",x"00",
-- [        ]
-- [   **   ]
-- [   **   ]
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"18",x"18",x"08",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [    *   ]
-- [        ]
x"00",x"00",x"00",x"3c",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [  ****  ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"02",x"06",x"0c",x"18",x"30",x"60",x"40",x"00",
-- [      * ]
-- [     ** ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ **     ]
-- [ *      ]
-- [        ]
x"3c",x"66",x"6e",x"7e",x"76",x"66",x"3c",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ ** *** ]
-- [ ****** ]
-- [ *** ** ]
-- [ **  ** ]
-- [  ****  ]
-- [        ]
x"18",x"38",x"18",x"18",x"18",x"18",x"7e",x"00",
-- [   **   ]
-- [  ***   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [ ****** ]
-- [        ]
x"7c",x"66",x"06",x"1c",x"30",x"66",x"7e",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [     ** ]
-- [   ***  ]
-- [  **    ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"7c",x"66",x"06",x"0c",x"06",x"66",x"7e",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [     ** ]
-- [    **  ]
-- [     ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"60",x"60",x"6c",x"7e",x"0c",x"0c",x"0c",x"00",
-- [ **     ]
-- [ **     ]
-- [ ** **  ]
-- [ ****** ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [        ]
x"7e",x"66",x"60",x"7c",x"06",x"66",x"7c",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [ **     ]
-- [ *****  ]
-- [     ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"3e",x"66",x"60",x"7c",x"66",x"66",x"3e",x"00",
-- [  ***** ]
-- [ **  ** ]
-- [ **     ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"7e",x"66",x"06",x"1e",x"06",x"06",x"06",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [     ** ]
-- [   **** ]
-- [     ** ]
-- [     ** ]
-- [     ** ]
-- [        ]
x"3c",x"66",x"66",x"3c",x"66",x"66",x"7e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"3c",x"66",x"66",x"3e",x"06",x"66",x"7c",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [     ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [        ]
x"00",x"18",x"18",x"00",x"18",x"18",x"08",x"00",
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [    *   ]
-- [        ]
x"00",x"0c",x"18",x"30",x"18",x"0c",x"00",x"00",
-- [        ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [   **   ]
-- [    **  ]
-- [        ]
-- [        ]
x"00",x"00",x"3c",x"00",x"3c",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [  ****  ]
-- [        ]
-- [  ****  ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"30",x"18",x"0c",x"18",x"30",x"00",x"00",
-- [        ]
-- [  **    ]
-- [   **   ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [        ]
-- [        ]
x"7e",x"66",x"06",x"0c",x"18",x"00",x"18",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [     ** ]
-- [    **  ]
-- [   **   ]
-- [        ]
-- [   **   ]
-- [        ]
x"00",x"00",x"00",x"ff",x"ff",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
x"08",x"1c",x"3e",x"7f",x"3e",x"1c",x"3e",x"00",
-- [    *   ]
-- [   ***  ]
-- [  ***** ]
-- [ *******]
-- [  ***** ]
-- [   ***  ]
-- [  ***** ]
-- [        ]
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"00",x"00",x"00",x"ff",x"ff",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"ff",x"ff",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",
-- [        ]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"ff",x"ff",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [        ]
-- [        ]
x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30",
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",x"0c",
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
x"00",x"00",x"00",x"e0",x"f0",x"38",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [***     ]
-- [****    ]
-- [  ***   ]
-- [   **   ]
-- [   **   ]
x"18",x"18",x"1c",x"0f",x"07",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   ***  ]
-- [    ****]
-- [     ***]
-- [        ]
-- [        ]
-- [        ]
x"18",x"18",x"38",x"f0",x"e0",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [  ***   ]
-- [****    ]
-- [***     ]
-- [        ]
-- [        ]
-- [        ]
x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"ff",x"ff",
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [********]
-- [********]
x"c0",x"e0",x"70",x"38",x"1c",x"0e",x"07",x"03",
-- [**      ]
-- [***     ]
-- [ ***    ]
-- [  ***   ]
-- [   ***  ]
-- [    *** ]
-- [     ***]
-- [      **]
x"03",x"07",x"0e",x"1c",x"38",x"70",x"e0",x"c0",
-- [      **]
-- [     ***]
-- [    *** ]
-- [   ***  ]
-- [  ***   ]
-- [ ***    ]
-- [***     ]
-- [**      ]
x"ff",x"ff",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",
-- [********]
-- [********]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
x"ff",x"ff",x"03",x"03",x"03",x"03",x"03",x"03",
-- [********]
-- [********]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
x"00",x"3c",x"7e",x"7e",x"7e",x"7e",x"3c",x"00",
-- [        ]
-- [  ****  ]
-- [ ****** ]
-- [ ****** ]
-- [ ****** ]
-- [ ****** ]
-- [  ****  ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [        ]
x"36",x"7f",x"7f",x"7f",x"3e",x"1c",x"08",x"00",
-- [  ** ** ]
-- [ *******]
-- [ *******]
-- [ *******]
-- [  ***** ]
-- [   ***  ]
-- [    *   ]
-- [        ]
x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
x"00",x"00",x"00",x"07",x"0f",x"1c",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [     ***]
-- [    ****]
-- [   ***  ]
-- [   **   ]
-- [   **   ]
x"c3",x"e7",x"7e",x"3c",x"3c",x"7e",x"e7",x"c3",
-- [**    **]
-- [***  ***]
-- [ ****** ]
-- [  ****  ]
-- [  ****  ]
-- [ ****** ]
-- [***  ***]
-- [**    **]
x"00",x"3c",x"66",x"42",x"42",x"66",x"3c",x"00",
-- [        ]
-- [  ****  ]
-- [ **  ** ]
-- [ *    * ]
-- [ *    * ]
-- [ **  ** ]
-- [  ****  ]
-- [        ]
x"18",x"18",x"7e",x"7e",x"18",x"18",x"3c",x"00",
-- [   **   ]
-- [   **   ]
-- [ ****** ]
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [  ****  ]
-- [        ]
x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",
-- [     ** ]
-- [     ** ]
-- [     ** ]
-- [     ** ]
-- [     ** ]
-- [     ** ]
-- [     ** ]
-- [     ** ]
x"08",x"1c",x"3e",x"7f",x"3e",x"1c",x"08",x"00",
-- [    *   ]
-- [   ***  ]
-- [  ***** ]
-- [ *******]
-- [  ***** ]
-- [   ***  ]
-- [    *   ]
-- [        ]
x"18",x"18",x"18",x"ff",x"ff",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [********]
-- [********]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"a0",x"50",x"a0",x"50",x"a0",x"50",x"a0",x"50",
-- [* *     ]
-- [ * *    ]
-- [* *     ]
-- [ * *    ]
-- [* *     ]
-- [ * *    ]
-- [* *     ]
-- [ * *    ]
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"00",x"00",x"00",x"3e",x"76",x"36",x"36",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [  ***** ]
-- [ *** ** ]
-- [  ** ** ]
-- [  ** ** ]
-- [        ]
x"ff",x"7f",x"3f",x"1f",x"0f",x"07",x"03",x"01",
-- [********]
-- [ *******]
-- [  ******]
-- [   *****]
-- [    ****]
-- [     ***]
-- [      **]
-- [       *]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
x"00",x"00",x"00",x"00",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
x"00",x"00",x"00",x"00",x"aa",x"55",x"aa",x"55",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
x"ff",x"fe",x"fc",x"f8",x"f0",x"e0",x"c0",x"80",
-- [********]
-- [******* ]
-- [******  ]
-- [*****   ]
-- [****    ]
-- [***     ]
-- [**      ]
-- [*       ]
x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
x"18",x"18",x"18",x"1f",x"1f",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   *****]
-- [   *****]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"00",x"00",x"00",x"00",x"0f",x"0f",x"0f",x"0f",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"18",x"18",x"18",x"1f",x"1f",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   *****]
-- [   *****]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"f8",x"f8",x"18",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [*****   ]
-- [*****   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
x"00",x"00",x"00",x"1f",x"1f",x"18",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [   *****]
-- [   *****]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"18",x"18",x"18",x"ff",x"ff",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"ff",x"ff",x"18",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"18",x"18",x"18",x"f8",x"f8",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [*****   ]
-- [*****   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
x"03",x"03",x"03",x"03",x"03",x"03",x"ff",x"ff",
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [********]
-- [********]
x"00",x"00",x"00",x"00",x"f0",x"f0",x"f0",x"f0",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
x"0f",x"0f",x"0f",x"0f",x"00",x"00",x"00",x"00",
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"18",x"18",x"18",x"f8",x"f8",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [*****   ]
-- [*****   ]
-- [        ]
-- [        ]
-- [        ]
x"f0",x"f0",x"f0",x"f0",x"00",x"00",x"00",x"00",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"f0",x"f0",x"f0",x"f0",x"0f",x"0f",x"0f",x"0f",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"c3",x"99",x"91",x"91",x"9f",x"99",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  *   *]
-- [*  *   *]
-- [*  *****]
-- [*  **  *]
-- [**     *]
-- [********]
x"c3",x"99",x"99",x"81",x"99",x"99",x"99",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"83",x"99",x"99",x"83",x"99",x"99",x"81",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"c3",x"99",x"99",x"9f",x"9f",x"99",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*  *****]
-- [*  *****]
-- [*  **  *]
-- [**     *]
-- [********]
x"83",x"99",x"99",x"99",x"99",x"99",x"83",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"81",x"99",x"9f",x"87",x"9f",x"99",x"81",x"ff",
-- [*      *]
-- [*  **  *]
-- [*  *****]
-- [*    ***]
-- [*  *****]
-- [*  **  *]
-- [*      *]
-- [********]
x"81",x"99",x"9f",x"87",x"9f",x"9f",x"9f",x"ff",
-- [*      *]
-- [*  **  *]
-- [*  *****]
-- [*    ***]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [********]
x"c1",x"99",x"9f",x"91",x"99",x"99",x"c1",x"ff",
-- [**     *]
-- [*  **  *]
-- [*  *****]
-- [*  *   *]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"99",x"99",x"99",x"81",x"99",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"81",x"e7",x"e7",x"e7",x"e7",x"e7",x"81",x"ff",
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [*      *]
-- [********]
x"81",x"99",x"f9",x"f9",x"99",x"99",x"83",x"ff",
-- [*      *]
-- [*  **  *]
-- [*****  *]
-- [*****  *]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"99",x"99",x"93",x"87",x"93",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  *  **]
-- [*    ***]
-- [*  *  **]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"9f",x"9f",x"9f",x"9f",x"9f",x"99",x"81",x"ff",
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  **  *]
-- [*      *]
-- [********]
x"9c",x"88",x"80",x"80",x"94",x"9c",x"9c",x"ff",
-- [*  ***  ]
-- [*   *   ]
-- [*       ]
-- [*       ]
-- [*  * *  ]
-- [*  ***  ]
-- [*  ***  ]
-- [********]
x"99",x"99",x"89",x"81",x"91",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*   *  *]
-- [*      *]
-- [*  *   *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"c3",x"99",x"99",x"99",x"99",x"99",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"83",x"99",x"99",x"81",x"9f",x"9f",x"9f",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [********]
x"c3",x"99",x"99",x"99",x"95",x"93",x"c9",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  * * *]
-- [*  *  **]
-- [**  *  *]
-- [********]
x"83",x"99",x"99",x"83",x"99",x"99",x"99",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"c1",x"9f",x"8f",x"c3",x"f1",x"f1",x"83",x"ff",
-- [**     *]
-- [*  *****]
-- [*   ****]
-- [**    **]
-- [****   *]
-- [****   *]
-- [*     **]
-- [********]
x"81",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"ff",
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [********]
x"99",x"99",x"99",x"99",x"99",x"91",x"c3",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  *   *]
-- [**    **]
-- [********]
x"99",x"99",x"99",x"d3",x"c3",x"e7",x"e7",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [** *  **]
-- [**    **]
-- [***  ***]
-- [***  ***]
-- [********]
x"9c",x"9c",x"94",x"80",x"80",x"88",x"9c",x"ff",
-- [*  ***  ]
-- [*  ***  ]
-- [*  * *  ]
-- [*       ]
-- [*       ]
-- [*   *   ]
-- [*  ***  ]
-- [********]
x"99",x"99",x"c3",x"e7",x"c3",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [**    **]
-- [***  ***]
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"99",x"99",x"91",x"c3",x"e7",x"e7",x"e7",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  *   *]
-- [**    **]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [********]
x"81",x"99",x"f3",x"e7",x"cf",x"89",x"81",x"ff",
-- [*      *]
-- [*  **  *]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [*   *  *]
-- [*      *]
-- [********]
x"c3",x"cf",x"cf",x"cf",x"cf",x"cf",x"c3",x"ff",
-- [**    **]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**    **]
-- [********]
x"c3",x"99",x"9f",x"87",x"cf",x"cf",x"81",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  *****]
-- [*    ***]
-- [**  ****]
-- [**  ****]
-- [*      *]
-- [********]
x"c3",x"f3",x"f3",x"f3",x"f3",x"f3",x"c3",x"ff",
-- [**    **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [**    **]
-- [********]
x"f7",x"e3",x"c1",x"e3",x"e3",x"e3",x"e3",x"ff",
-- [**** ***]
-- [***   **]
-- [**     *]
-- [***   **]
-- [***   **]
-- [***   **]
-- [***   **]
-- [********]
x"ff",x"ef",x"c0",x"80",x"c0",x"ef",x"ff",x"ff",
-- [********]
-- [*** ****]
-- [**      ]
-- [*       ]
-- [**      ]
-- [*** ****]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"c7",x"c7",x"c7",x"c7",x"c7",x"ff",x"c7",x"ff",
-- [**   ***]
-- [**   ***]
-- [**   ***]
-- [**   ***]
-- [**   ***]
-- [********]
-- [**   ***]
-- [********]
x"93",x"93",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [*  *  **]
-- [*  *  **]
-- [* ** ***]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"c9",x"c9",x"80",x"c9",x"80",x"c9",x"c9",x"ff",
-- [**  *  *]
-- [**  *  *]
-- [*       ]
-- [**  *  *]
-- [*       ]
-- [**  *  *]
-- [**  *  *]
-- [********]
x"e7",x"81",x"9f",x"81",x"f9",x"81",x"e7",x"ff",
-- [***  ***]
-- [*      *]
-- [*  *****]
-- [*      *]
-- [*****  *]
-- [*      *]
-- [***  ***]
-- [********]
x"9d",x"99",x"f3",x"e7",x"cf",x"99",x"b9",x"ff",
-- [*  *** *]
-- [*  **  *]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [*  **  *]
-- [* ***  *]
-- [********]
x"c3",x"99",x"99",x"c3",x"8b",x"91",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [**    **]
-- [*   * **]
-- [*  *   *]
-- [**     *]
-- [********]
x"e7",x"e7",x"ef",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [*** ****]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"e3",x"cf",x"cf",x"cf",x"cf",x"cf",x"e3",x"ff",
-- [***   **]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [***   **]
-- [********]
x"c7",x"f3",x"f3",x"f3",x"f3",x"f3",x"c7",x"ff",
-- [**   ***]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [**   ***]
-- [********]
x"f7",x"d5",x"e3",x"80",x"e3",x"d5",x"f7",x"ff",
-- [**** ***]
-- [** * * *]
-- [***   **]
-- [*       ]
-- [***   **]
-- [** * * *]
-- [**** ***]
-- [********]
x"ff",x"e7",x"e7",x"81",x"e7",x"e7",x"ff",x"ff",
-- [********]
-- [***  ***]
-- [***  ***]
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"e7",x"e7",x"f7",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [***  ***]
-- [***  ***]
-- [**** ***]
-- [********]
x"ff",x"ff",x"ff",x"c3",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [**    **]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"e7",x"e7",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
x"fd",x"f9",x"f3",x"e7",x"cf",x"9f",x"bf",x"ff",
-- [****** *]
-- [*****  *]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [*  *****]
-- [* ******]
-- [********]
x"c3",x"99",x"91",x"81",x"89",x"99",x"c3",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  *   *]
-- [*      *]
-- [*   *  *]
-- [*  **  *]
-- [**    **]
-- [********]
x"e7",x"c7",x"e7",x"e7",x"e7",x"e7",x"81",x"ff",
-- [***  ***]
-- [**   ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [*      *]
-- [********]
x"83",x"99",x"f9",x"e3",x"cf",x"99",x"81",x"ff",
-- [*     **]
-- [*  **  *]
-- [*****  *]
-- [***   **]
-- [**  ****]
-- [*  **  *]
-- [*      *]
-- [********]
x"83",x"99",x"f9",x"f3",x"f9",x"99",x"81",x"ff",
-- [*     **]
-- [*  **  *]
-- [*****  *]
-- [****  **]
-- [*****  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"9f",x"9f",x"93",x"81",x"f3",x"f3",x"f3",x"ff",
-- [*  *****]
-- [*  *****]
-- [*  *  **]
-- [*      *]
-- [****  **]
-- [****  **]
-- [****  **]
-- [********]
x"81",x"99",x"9f",x"83",x"f9",x"99",x"83",x"ff",
-- [*      *]
-- [*  **  *]
-- [*  *****]
-- [*     **]
-- [*****  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"c1",x"99",x"9f",x"83",x"99",x"99",x"c1",x"ff",
-- [**     *]
-- [*  **  *]
-- [*  *****]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"81",x"99",x"f9",x"e1",x"f9",x"f9",x"f9",x"ff",
-- [*      *]
-- [*  **  *]
-- [*****  *]
-- [***    *]
-- [*****  *]
-- [*****  *]
-- [*****  *]
-- [********]
x"c3",x"99",x"99",x"c3",x"99",x"99",x"81",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"c3",x"99",x"99",x"c1",x"f9",x"99",x"83",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [*****  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"ff",x"e7",x"e7",x"ff",x"e7",x"e7",x"ff",x"ff",
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
-- [********]
x"ff",x"e7",x"e7",x"ff",x"e7",x"e7",x"f7",x"ff",
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
-- [***  ***]
-- [***  ***]
-- [**** ***]
-- [********]
x"ff",x"f3",x"e7",x"cf",x"e7",x"f3",x"ff",x"ff",
-- [********]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [***  ***]
-- [****  **]
-- [********]
-- [********]
x"ff",x"ff",x"c3",x"ff",x"c3",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [**    **]
-- [********]
-- [**    **]
-- [********]
-- [********]
-- [********]
x"ff",x"cf",x"e7",x"f3",x"e7",x"cf",x"ff",x"ff",
-- [********]
-- [**  ****]
-- [***  ***]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [********]
-- [********]
x"81",x"99",x"f9",x"f3",x"e7",x"ff",x"e7",x"ff",
-- [*      *]
-- [*  **  *]
-- [*****  *]
-- [****  **]
-- [***  ***]
-- [********]
-- [***  ***]
-- [********]
x"ff",x"ff",x"ff",x"00",x"00",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
x"f7",x"e3",x"c1",x"80",x"c1",x"e3",x"c1",x"ff",
-- [**** ***]
-- [***   **]
-- [**     *]
-- [*       ]
-- [**     *]
-- [***   **]
-- [**     *]
-- [********]
x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"ff",x"ff",x"ff",x"00",x"00",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"00",x"00",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [********]
-- [********]
x"cf",x"cf",x"cf",x"cf",x"cf",x"cf",x"cf",x"cf",
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
x"f3",x"f3",x"f3",x"f3",x"f3",x"f3",x"f3",x"f3",
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
x"ff",x"ff",x"ff",x"1f",x"0f",x"c7",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [   *****]
-- [    ****]
-- [**   ***]
-- [***  ***]
-- [***  ***]
x"e7",x"e7",x"e3",x"f0",x"f8",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [***   **]
-- [****    ]
-- [*****   ]
-- [********]
-- [********]
-- [********]
x"e7",x"e7",x"c7",x"0f",x"1f",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [**   ***]
-- [    ****]
-- [   *****]
-- [********]
-- [********]
-- [********]
x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"00",x"00",
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [        ]
-- [        ]
x"3f",x"1f",x"8f",x"c7",x"e3",x"f1",x"f8",x"fc",
-- [  ******]
-- [   *****]
-- [*   ****]
-- [**   ***]
-- [***   **]
-- [****   *]
-- [*****   ]
-- [******  ]
x"fc",x"f8",x"f1",x"e3",x"c7",x"8f",x"1f",x"3f",
-- [******  ]
-- [*****   ]
-- [****   *]
-- [***   **]
-- [**   ***]
-- [*   ****]
-- [   *****]
-- [  ******]
x"00",x"00",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",
-- [        ]
-- [        ]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
x"00",x"00",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",
-- [        ]
-- [        ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
x"ff",x"c3",x"81",x"81",x"81",x"81",x"c3",x"ff",
-- [********]
-- [**    **]
-- [*      *]
-- [*      *]
-- [*      *]
-- [*      *]
-- [**    **]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [********]
x"c9",x"80",x"80",x"80",x"c1",x"e3",x"f7",x"ff",
-- [**  *  *]
-- [*       ]
-- [*       ]
-- [*       ]
-- [**     *]
-- [***   **]
-- [**** ***]
-- [********]
x"9f",x"9f",x"9f",x"9f",x"9f",x"9f",x"9f",x"9f",
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
x"ff",x"ff",x"ff",x"f8",x"f0",x"e3",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [*****   ]
-- [****    ]
-- [***   **]
-- [***  ***]
-- [***  ***]
x"3c",x"18",x"81",x"c3",x"c3",x"81",x"18",x"3c",
-- [  ****  ]
-- [   **   ]
-- [*      *]
-- [**    **]
-- [**    **]
-- [*      *]
-- [   **   ]
-- [  ****  ]
x"ff",x"c3",x"99",x"bd",x"bd",x"99",x"c3",x"ff",
-- [********]
-- [**    **]
-- [*  **  *]
-- [* **** *]
-- [* **** *]
-- [*  **  *]
-- [**    **]
-- [********]
x"e7",x"e7",x"81",x"81",x"e7",x"e7",x"c3",x"ff",
-- [***  ***]
-- [***  ***]
-- [*      *]
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [**    **]
-- [********]
x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",
-- [*****  *]
-- [*****  *]
-- [*****  *]
-- [*****  *]
-- [*****  *]
-- [*****  *]
-- [*****  *]
-- [*****  *]
x"f7",x"e3",x"c1",x"80",x"c1",x"e3",x"f7",x"ff",
-- [**** ***]
-- [***   **]
-- [**     *]
-- [*       ]
-- [**     *]
-- [***   **]
-- [**** ***]
-- [********]
x"e7",x"e7",x"e7",x"00",x"00",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [        ]
-- [        ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"5f",x"af",x"5f",x"af",x"5f",x"af",x"5f",x"af",
-- [ * *****]
-- [* * ****]
-- [ * *****]
-- [* * ****]
-- [ * *****]
-- [* * ****]
-- [ * *****]
-- [* * ****]
x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"ff",x"ff",x"ff",x"c1",x"89",x"c9",x"c9",x"ff",
-- [********]
-- [********]
-- [********]
-- [**     *]
-- [*   *  *]
-- [**  *  *]
-- [**  *  *]
-- [********]
x"00",x"80",x"c0",x"e0",x"f0",x"f8",x"fc",x"fe",
-- [        ]
-- [*       ]
-- [**      ]
-- [***     ]
-- [****    ]
-- [*****   ]
-- [******  ]
-- [******* ]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
x"ff",x"ff",x"ff",x"ff",x"55",x"aa",x"55",x"aa",
-- [********]
-- [********]
-- [********]
-- [********]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
x"00",x"01",x"03",x"07",x"0f",x"1f",x"3f",x"7f",
-- [        ]
-- [       *]
-- [      **]
-- [     ***]
-- [    ****]
-- [   *****]
-- [  ******]
-- [ *******]
x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
x"e7",x"e7",x"e7",x"e0",x"e0",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***     ]
-- [***     ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"ff",x"ff",x"ff",x"ff",x"f0",x"f0",x"f0",x"f0",
-- [********]
-- [********]
-- [********]
-- [********]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
x"e7",x"e7",x"e7",x"e0",x"e0",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***     ]
-- [***     ]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"07",x"07",x"e7",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [     ***]
-- [     ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
x"ff",x"ff",x"ff",x"e0",x"e0",x"e7",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [***     ]
-- [***     ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"e7",x"e7",x"e7",x"00",x"00",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"00",x"00",x"e7",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"e7",x"e7",x"e7",x"07",x"07",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [     ***]
-- [     ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
x"1f",x"1f",x"1f",x"1f",x"1f",x"1f",x"1f",x"1f",
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"00",x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"00",x"00",
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [        ]
-- [        ]
x"ff",x"ff",x"ff",x"ff",x"0f",x"0f",x"0f",x"0f",
-- [********]
-- [********]
-- [********]
-- [********]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"f0",x"f0",x"f0",x"f0",x"ff",x"ff",x"ff",x"ff",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [********]
-- [********]
-- [********]
-- [********]
x"e7",x"e7",x"e7",x"07",x"07",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [     ***]
-- [     ***]
-- [********]
-- [********]
-- [********]
x"0f",x"0f",x"0f",x"0f",x"ff",x"ff",x"ff",x"ff",
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [********]
-- [********]
-- [********]
-- [********]
x"0f",x"0f",x"0f",x"0f",x"f0",x"f0",x"f0",x"f0",
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
x"3c",x"66",x"6e",x"6e",x"60",x"66",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ ** *** ]
-- [ ** *** ]
-- [ **     ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"00",x"00",x"3c",x"06",x"3e",x"66",x"7e",x"00",
-- [        ]
-- [        ]
-- [  ****  ]
-- [     ** ]
-- [  ***** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"00",x"60",x"60",x"7c",x"66",x"66",x"7e",x"00",
-- [        ]
-- [ **     ]
-- [ **     ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"00",x"00",x"3e",x"60",x"60",x"60",x"7e",x"00",
-- [        ]
-- [        ]
-- [  ***** ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ ****** ]
-- [        ]
x"00",x"06",x"06",x"3e",x"66",x"66",x"7e",x"00",
-- [        ]
-- [     ** ]
-- [     ** ]
-- [  ***** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"00",x"00",x"3c",x"66",x"7e",x"60",x"7e",x"00",
-- [        ]
-- [        ]
-- [  ****  ]
-- [ **  ** ]
-- [ ****** ]
-- [ **     ]
-- [ ****** ]
-- [        ]
x"00",x"0e",x"18",x"3c",x"18",x"18",x"18",x"00",
-- [        ]
-- [    *** ]
-- [   **   ]
-- [  ****  ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"00",x"00",x"3e",x"66",x"66",x"7e",x"06",x"3c",
-- [        ]
-- [        ]
-- [  ***** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [     ** ]
-- [  ****  ]
x"00",x"60",x"60",x"7c",x"66",x"66",x"66",x"00",
-- [        ]
-- [ **     ]
-- [ **     ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"00",x"18",x"00",x"18",x"18",x"18",x"18",x"00",
-- [        ]
-- [   **   ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"00",x"0c",x"00",x"0c",x"0c",x"0c",x"6c",x"78",
-- [        ]
-- [    **  ]
-- [        ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [ ** **  ]
-- [ ****   ]
x"00",x"60",x"66",x"6c",x"78",x"6c",x"66",x"00",
-- [        ]
-- [ **     ]
-- [ **  ** ]
-- [ ** **  ]
-- [ ****   ]
-- [ ** **  ]
-- [ **  ** ]
-- [        ]
x"00",x"18",x"18",x"18",x"18",x"18",x"3c",x"00",
-- [        ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [  ****  ]
-- [        ]
x"00",x"00",x"7e",x"6b",x"6b",x"63",x"63",x"00",
-- [        ]
-- [        ]
-- [ ****** ]
-- [ ** * **]
-- [ ** * **]
-- [ **   **]
-- [ **   **]
-- [        ]
x"00",x"00",x"7c",x"66",x"66",x"66",x"66",x"00",
-- [        ]
-- [        ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"00",x"00",x"3c",x"66",x"66",x"66",x"3e",x"00",
-- [        ]
-- [        ]
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"00",x"00",x"7c",x"66",x"66",x"7e",x"60",x"60",
-- [        ]
-- [        ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [ **     ]
-- [ **     ]
x"00",x"00",x"3e",x"66",x"66",x"7e",x"06",x"06",
-- [        ]
-- [        ]
-- [  ***** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [     ** ]
-- [     ** ]
x"00",x"00",x"7e",x"66",x"60",x"60",x"60",x"00",
-- [        ]
-- [        ]
-- [ ****** ]
-- [ **  ** ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [        ]
x"00",x"00",x"3e",x"60",x"7e",x"06",x"7e",x"00",
-- [        ]
-- [        ]
-- [  ***** ]
-- [ **     ]
-- [ ****** ]
-- [     ** ]
-- [ ****** ]
-- [        ]
x"00",x"18",x"7e",x"18",x"18",x"18",x"1c",x"00",
-- [        ]
-- [   **   ]
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   ***  ]
-- [        ]
x"00",x"00",x"66",x"66",x"66",x"66",x"3e",x"00",
-- [        ]
-- [        ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"00",x"00",x"66",x"66",x"66",x"34",x"18",x"00",
-- [        ]
-- [        ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ** *  ]
-- [   **   ]
-- [        ]
x"00",x"00",x"63",x"63",x"6b",x"6b",x"3f",x"00",
-- [        ]
-- [        ]
-- [ **   **]
-- [ **   **]
-- [ ** * **]
-- [ ** * **]
-- [  ******]
-- [        ]
x"00",x"00",x"66",x"3c",x"18",x"3c",x"66",x"00",
-- [        ]
-- [        ]
-- [ **  ** ]
-- [  ****  ]
-- [   **   ]
-- [  ****  ]
-- [ **  ** ]
-- [        ]
x"00",x"00",x"66",x"66",x"66",x"3c",x"18",x"30",
-- [        ]
-- [        ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ****  ]
-- [   **   ]
-- [  **    ]
x"00",x"00",x"7e",x"0c",x"18",x"30",x"7e",x"00",
-- [        ]
-- [        ]
-- [ ****** ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ ****** ]
-- [        ]
x"3c",x"30",x"30",x"30",x"30",x"30",x"3c",x"00",
-- [  ****  ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  ****  ]
-- [        ]
x"3c",x"66",x"60",x"78",x"30",x"30",x"7e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **     ]
-- [ ****   ]
-- [  **    ]
-- [  **    ]
-- [ ****** ]
-- [        ]
x"3c",x"0c",x"0c",x"0c",x"0c",x"0c",x"3c",x"00",
-- [  ****  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [  ****  ]
-- [        ]
x"08",x"1c",x"3e",x"1c",x"1c",x"1c",x"1c",x"00",
-- [    *   ]
-- [   ***  ]
-- [  ***** ]
-- [   ***  ]
-- [   ***  ]
-- [   ***  ]
-- [   ***  ]
-- [        ]
x"00",x"10",x"3f",x"7f",x"3f",x"10",x"00",x"00",
-- [        ]
-- [   *    ]
-- [  ******]
-- [ *******]
-- [  ******]
-- [   *    ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"38",x"38",x"38",x"38",x"38",x"00",x"38",x"00",
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [  ***   ]
-- [        ]
-- [  ***   ]
-- [        ]
x"6c",x"6c",x"48",x"00",x"00",x"00",x"00",x"00",
-- [ ** **  ]
-- [ ** **  ]
-- [ *  *   ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"36",x"36",x"7f",x"36",x"7f",x"36",x"36",x"00",
-- [  ** ** ]
-- [  ** ** ]
-- [ *******]
-- [  ** ** ]
-- [ *******]
-- [  ** ** ]
-- [  ** ** ]
-- [        ]
x"18",x"7e",x"60",x"7e",x"06",x"7e",x"18",x"00",
-- [   **   ]
-- [ ****** ]
-- [ **     ]
-- [ ****** ]
-- [     ** ]
-- [ ****** ]
-- [   **   ]
-- [        ]
x"62",x"66",x"0c",x"18",x"30",x"66",x"46",x"00",
-- [ **   * ]
-- [ **  ** ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ **  ** ]
-- [ *   ** ]
-- [        ]
x"3c",x"66",x"66",x"3c",x"74",x"6e",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ****  ]
-- [ *** *  ]
-- [ ** *** ]
-- [  ***** ]
-- [        ]
x"18",x"18",x"10",x"00",x"00",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   *    ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"1c",x"30",x"30",x"30",x"30",x"30",x"1c",x"00",
-- [   ***  ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [  **    ]
-- [   ***  ]
-- [        ]
x"38",x"0c",x"0c",x"0c",x"0c",x"0c",x"38",x"00",
-- [  ***   ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [  ***   ]
-- [        ]
x"08",x"2a",x"1c",x"7f",x"1c",x"2a",x"08",x"00",
-- [    *   ]
-- [  * * * ]
-- [   ***  ]
-- [ *******]
-- [   ***  ]
-- [  * * * ]
-- [    *   ]
-- [        ]
x"00",x"18",x"18",x"7e",x"18",x"18",x"00",x"00",
-- [        ]
-- [   **   ]
-- [   **   ]
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"18",x"18",x"08",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [    *   ]
-- [        ]
x"00",x"00",x"00",x"3c",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [  ****  ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"02",x"06",x"0c",x"18",x"30",x"60",x"40",x"00",
-- [      * ]
-- [     ** ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ **     ]
-- [ *      ]
-- [        ]
x"3c",x"66",x"6e",x"7e",x"76",x"66",x"3c",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ ** *** ]
-- [ ****** ]
-- [ *** ** ]
-- [ **  ** ]
-- [  ****  ]
-- [        ]
x"18",x"38",x"18",x"18",x"18",x"18",x"7e",x"00",
-- [   **   ]
-- [  ***   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [ ****** ]
-- [        ]
x"7c",x"66",x"06",x"1c",x"30",x"66",x"7e",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [     ** ]
-- [   ***  ]
-- [  **    ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"7c",x"66",x"06",x"0c",x"06",x"66",x"7e",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [     ** ]
-- [    **  ]
-- [     ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"60",x"60",x"6c",x"7e",x"0c",x"0c",x"0c",x"00",
-- [ **     ]
-- [ **     ]
-- [ ** **  ]
-- [ ****** ]
-- [    **  ]
-- [    **  ]
-- [    **  ]
-- [        ]
x"7e",x"66",x"60",x"7c",x"06",x"66",x"7c",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [ **     ]
-- [ *****  ]
-- [     ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"3e",x"66",x"60",x"7c",x"66",x"66",x"3e",x"00",
-- [  ***** ]
-- [ **  ** ]
-- [ **     ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"7e",x"66",x"06",x"1e",x"06",x"06",x"06",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [     ** ]
-- [   **** ]
-- [     ** ]
-- [     ** ]
-- [     ** ]
-- [        ]
x"3c",x"66",x"66",x"3c",x"66",x"66",x"7e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"3c",x"66",x"66",x"3e",x"06",x"66",x"7c",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [     ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"00",x"18",x"18",x"00",x"18",x"18",x"00",x"00",
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [        ]
x"00",x"18",x"18",x"00",x"18",x"18",x"08",x"00",
-- [        ]
-- [   **   ]
-- [   **   ]
-- [        ]
-- [   **   ]
-- [   **   ]
-- [    *   ]
-- [        ]
x"00",x"0c",x"18",x"30",x"18",x"0c",x"00",x"00",
-- [        ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [   **   ]
-- [    **  ]
-- [        ]
-- [        ]
x"00",x"00",x"3c",x"00",x"3c",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [  ****  ]
-- [        ]
-- [  ****  ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"30",x"18",x"0c",x"18",x"30",x"00",x"00",
-- [        ]
-- [  **    ]
-- [   **   ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [        ]
-- [        ]
x"7e",x"66",x"06",x"0c",x"18",x"00",x"18",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [     ** ]
-- [    **  ]
-- [   **   ]
-- [        ]
-- [   **   ]
-- [        ]
x"00",x"00",x"00",x"ff",x"ff",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
x"3c",x"66",x"66",x"7e",x"66",x"66",x"66",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"7c",x"66",x"66",x"7c",x"66",x"66",x"7e",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"3c",x"66",x"66",x"60",x"60",x"66",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **     ]
-- [ **     ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"7c",x"66",x"66",x"66",x"66",x"66",x"7c",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"7e",x"66",x"60",x"78",x"60",x"66",x"7e",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [ **     ]
-- [ ****   ]
-- [ **     ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"7e",x"66",x"60",x"78",x"60",x"60",x"60",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [ **     ]
-- [ ****   ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [        ]
x"3e",x"66",x"60",x"6e",x"66",x"66",x"3e",x"00",
-- [  ***** ]
-- [ **  ** ]
-- [ **     ]
-- [ ** *** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"66",x"66",x"66",x"7e",x"66",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"7e",x"18",x"18",x"18",x"18",x"18",x"7e",x"00",
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [ ****** ]
-- [        ]
x"7e",x"66",x"06",x"06",x"66",x"66",x"7c",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [     ** ]
-- [     ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [        ]
x"66",x"66",x"6c",x"78",x"6c",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ ** **  ]
-- [ ****   ]
-- [ ** **  ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"60",x"60",x"60",x"60",x"60",x"66",x"7e",x"00",
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [ **  ** ]
-- [ ****** ]
-- [        ]
x"63",x"77",x"7f",x"7f",x"6b",x"63",x"63",x"00",
-- [ **   **]
-- [ *** ***]
-- [ *******]
-- [ *******]
-- [ ** * **]
-- [ **   **]
-- [ **   **]
-- [        ]
x"66",x"66",x"76",x"7e",x"6e",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ *** ** ]
-- [ ****** ]
-- [ ** *** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"3c",x"66",x"66",x"66",x"66",x"66",x"3e",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  ***** ]
-- [        ]
x"7c",x"66",x"66",x"7e",x"60",x"60",x"60",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ****** ]
-- [ **     ]
-- [ **     ]
-- [ **     ]
-- [        ]
x"3c",x"66",x"66",x"66",x"6a",x"6c",x"36",x"00",
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ** * * ]
-- [ ** **  ]
-- [  ** ** ]
-- [        ]
x"7c",x"66",x"66",x"7c",x"66",x"66",x"66",x"00",
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ *****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"3e",x"60",x"70",x"3c",x"0e",x"0e",x"7c",x"00",
-- [  ***** ]
-- [ **     ]
-- [ ***    ]
-- [  ****  ]
-- [    *** ]
-- [    *** ]
-- [ *****  ]
-- [        ]
x"7e",x"18",x"18",x"18",x"18",x"18",x"18",x"00",
-- [ ****** ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"66",x"66",x"66",x"66",x"66",x"6e",x"3c",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [ ** *** ]
-- [  ****  ]
-- [        ]
x"66",x"66",x"66",x"2c",x"3c",x"18",x"18",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ **  ** ]
-- [  * **  ]
-- [  ****  ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"63",x"63",x"6b",x"7f",x"7f",x"77",x"63",x"00",
-- [ **   **]
-- [ **   **]
-- [ ** * **]
-- [ *******]
-- [ *******]
-- [ *** ***]
-- [ **   **]
-- [        ]
x"66",x"66",x"3c",x"18",x"3c",x"66",x"66",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [  ****  ]
-- [   **   ]
-- [  ****  ]
-- [ **  ** ]
-- [ **  ** ]
-- [        ]
x"66",x"66",x"6e",x"3c",x"18",x"18",x"18",x"00",
-- [ **  ** ]
-- [ **  ** ]
-- [ ** *** ]
-- [  ****  ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [        ]
x"7e",x"66",x"0c",x"18",x"30",x"76",x"7e",x"00",
-- [ ****** ]
-- [ **  ** ]
-- [    **  ]
-- [   **   ]
-- [  **    ]
-- [ *** ** ]
-- [ ****** ]
-- [        ]
x"18",x"18",x"18",x"ff",x"ff",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [********]
-- [********]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"c0",x"c0",x"30",x"30",x"c0",x"c0",x"30",x"30",
-- [**      ]
-- [**      ]
-- [  **    ]
-- [  **    ]
-- [**      ]
-- [**      ]
-- [  **    ]
-- [  **    ]
x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
x"33",x"99",x"cc",x"66",x"33",x"99",x"cc",x"66",
-- [  **  **]
-- [*  **  *]
-- [**  **  ]
-- [ **  ** ]
-- [  **  **]
-- [*  **  *]
-- [**  **  ]
-- [ **  ** ]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
x"00",x"00",x"00",x"00",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
x"00",x"00",x"00",x"00",x"aa",x"55",x"aa",x"55",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
x"cc",x"99",x"33",x"66",x"cc",x"99",x"33",x"66",
-- [**  **  ]
-- [*  **  *]
-- [  **  **]
-- [ **  ** ]
-- [**  **  ]
-- [*  **  *]
-- [  **  **]
-- [ **  ** ]
x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
-- [      **]
x"18",x"18",x"18",x"1f",x"1f",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   *****]
-- [   *****]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"00",x"00",x"00",x"00",x"0f",x"0f",x"0f",x"0f",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"18",x"18",x"18",x"1f",x"1f",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [   *****]
-- [   *****]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"f8",x"f8",x"18",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [*****   ]
-- [*****   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"00",x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
x"00",x"00",x"00",x"1f",x"1f",x"18",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [   *****]
-- [   *****]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"18",x"18",x"18",x"ff",x"ff",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"ff",x"ff",x"18",x"18",x"18",
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"18",x"18",x"18",x"f8",x"f8",x"18",x"18",x"18",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [*****   ]
-- [*****   ]
-- [   **   ]
-- [   **   ]
-- [   **   ]
x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
-- [**      ]
x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
-- [***     ]
x"07",x"07",x"07",x"07",x"07",x"07",x"07",x"07",
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
-- [     ***]
x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",x"00",
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"00",x"00",x"00",x"00",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
x"00",x"01",x"03",x"46",x"6c",x"38",x"10",x"00",
-- [        ]
-- [       *]
-- [      **]
-- [ *   ** ]
-- [ ** **  ]
-- [  ***   ]
-- [   *    ]
-- [        ]
x"00",x"00",x"00",x"00",x"f0",x"f0",x"f0",x"f0",
-- [        ]
-- [        ]
-- [        ]
-- [        ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
x"0f",x"0f",x"0f",x"0f",x"00",x"00",x"00",x"00",
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"18",x"18",x"18",x"f8",x"f8",x"00",x"00",x"00",
-- [   **   ]
-- [   **   ]
-- [   **   ]
-- [*****   ]
-- [*****   ]
-- [        ]
-- [        ]
-- [        ]
x"f0",x"f0",x"f0",x"f0",x"00",x"00",x"00",x"00",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"f0",x"f0",x"f0",x"f0",x"0f",x"0f",x"0f",x"0f",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"c3",x"99",x"91",x"91",x"9f",x"99",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  *   *]
-- [*  *   *]
-- [*  *****]
-- [*  **  *]
-- [**     *]
-- [********]
x"ff",x"ff",x"c3",x"f9",x"c1",x"99",x"81",x"ff",
-- [********]
-- [********]
-- [**    **]
-- [*****  *]
-- [**     *]
-- [*  **  *]
-- [*      *]
-- [********]
x"ff",x"9f",x"9f",x"83",x"99",x"99",x"81",x"ff",
-- [********]
-- [*  *****]
-- [*  *****]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"ff",x"ff",x"c1",x"9f",x"9f",x"9f",x"81",x"ff",
-- [********]
-- [********]
-- [**     *]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*      *]
-- [********]
x"ff",x"f9",x"f9",x"c1",x"99",x"99",x"81",x"ff",
-- [********]
-- [*****  *]
-- [*****  *]
-- [**     *]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"ff",x"ff",x"c3",x"99",x"81",x"9f",x"81",x"ff",
-- [********]
-- [********]
-- [**    **]
-- [*  **  *]
-- [*      *]
-- [*  *****]
-- [*      *]
-- [********]
x"ff",x"f1",x"e7",x"c3",x"e7",x"e7",x"e7",x"ff",
-- [********]
-- [****   *]
-- [***  ***]
-- [**    **]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [********]
x"ff",x"ff",x"c1",x"99",x"99",x"81",x"f9",x"c3",
-- [********]
-- [********]
-- [**     *]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*****  *]
-- [**    **]
x"ff",x"9f",x"9f",x"83",x"99",x"99",x"99",x"ff",
-- [********]
-- [*  *****]
-- [*  *****]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"ff",x"e7",x"ff",x"e7",x"e7",x"e7",x"e7",x"ff",
-- [********]
-- [***  ***]
-- [********]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [********]
x"ff",x"f3",x"ff",x"f3",x"f3",x"f3",x"93",x"87",
-- [********]
-- [****  **]
-- [********]
-- [****  **]
-- [****  **]
-- [****  **]
-- [*  *  **]
-- [*    ***]
x"ff",x"9f",x"99",x"93",x"87",x"93",x"99",x"ff",
-- [********]
-- [*  *****]
-- [*  **  *]
-- [*  *  **]
-- [*    ***]
-- [*  *  **]
-- [*  **  *]
-- [********]
x"ff",x"e7",x"e7",x"e7",x"e7",x"e7",x"c3",x"ff",
-- [********]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [**    **]
-- [********]
x"ff",x"ff",x"81",x"94",x"94",x"9c",x"9c",x"ff",
-- [********]
-- [********]
-- [*      *]
-- [*  * *  ]
-- [*  * *  ]
-- [*  ***  ]
-- [*  ***  ]
-- [********]
x"ff",x"ff",x"83",x"99",x"99",x"99",x"99",x"ff",
-- [********]
-- [********]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"ff",x"ff",x"c3",x"99",x"99",x"99",x"c1",x"ff",
-- [********]
-- [********]
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"ff",x"ff",x"83",x"99",x"99",x"81",x"9f",x"9f",
-- [********]
-- [********]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*  *****]
-- [*  *****]
x"ff",x"ff",x"c1",x"99",x"99",x"81",x"f9",x"f9",
-- [********]
-- [********]
-- [**     *]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*****  *]
-- [*****  *]
x"ff",x"ff",x"81",x"99",x"9f",x"9f",x"9f",x"ff",
-- [********]
-- [********]
-- [*      *]
-- [*  **  *]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [********]
x"ff",x"ff",x"c1",x"9f",x"81",x"f9",x"81",x"ff",
-- [********]
-- [********]
-- [**     *]
-- [*  *****]
-- [*      *]
-- [*****  *]
-- [*      *]
-- [********]
x"ff",x"e7",x"81",x"e7",x"e7",x"e7",x"e3",x"ff",
-- [********]
-- [***  ***]
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***   **]
-- [********]
x"ff",x"ff",x"99",x"99",x"99",x"99",x"c1",x"ff",
-- [********]
-- [********]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"ff",x"ff",x"99",x"99",x"99",x"cb",x"e7",x"ff",
-- [********]
-- [********]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [**  * **]
-- [***  ***]
-- [********]
x"ff",x"ff",x"9c",x"9c",x"94",x"94",x"c0",x"ff",
-- [********]
-- [********]
-- [*  ***  ]
-- [*  ***  ]
-- [*  * *  ]
-- [*  * *  ]
-- [**      ]
-- [********]
x"ff",x"ff",x"99",x"c3",x"e7",x"c3",x"99",x"ff",
-- [********]
-- [********]
-- [*  **  *]
-- [**    **]
-- [***  ***]
-- [**    **]
-- [*  **  *]
-- [********]
x"ff",x"ff",x"99",x"99",x"99",x"c3",x"e7",x"cf",
-- [********]
-- [********]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [**    **]
-- [***  ***]
-- [**  ****]
x"ff",x"ff",x"81",x"f3",x"e7",x"cf",x"81",x"ff",
-- [********]
-- [********]
-- [*      *]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [*      *]
-- [********]
x"c3",x"cf",x"cf",x"cf",x"cf",x"cf",x"c3",x"ff",
-- [**    **]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**    **]
-- [********]
x"c3",x"99",x"9f",x"87",x"cf",x"cf",x"81",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  *****]
-- [*    ***]
-- [**  ****]
-- [**  ****]
-- [*      *]
-- [********]
x"c3",x"f3",x"f3",x"f3",x"f3",x"f3",x"c3",x"ff",
-- [**    **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [**    **]
-- [********]
x"f7",x"e3",x"c1",x"e3",x"e3",x"e3",x"e3",x"ff",
-- [**** ***]
-- [***   **]
-- [**     *]
-- [***   **]
-- [***   **]
-- [***   **]
-- [***   **]
-- [********]
x"ff",x"ef",x"c0",x"80",x"c0",x"ef",x"ff",x"ff",
-- [********]
-- [*** ****]
-- [**      ]
-- [*       ]
-- [**      ]
-- [*** ****]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"c7",x"c7",x"c7",x"c7",x"c7",x"ff",x"c7",x"ff",
-- [**   ***]
-- [**   ***]
-- [**   ***]
-- [**   ***]
-- [**   ***]
-- [********]
-- [**   ***]
-- [********]
x"93",x"93",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [*  *  **]
-- [*  *  **]
-- [* ** ***]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"c9",x"c9",x"80",x"c9",x"80",x"c9",x"c9",x"ff",
-- [**  *  *]
-- [**  *  *]
-- [*       ]
-- [**  *  *]
-- [*       ]
-- [**  *  *]
-- [**  *  *]
-- [********]
x"e7",x"81",x"9f",x"81",x"f9",x"81",x"e7",x"ff",
-- [***  ***]
-- [*      *]
-- [*  *****]
-- [*      *]
-- [*****  *]
-- [*      *]
-- [***  ***]
-- [********]
x"9d",x"99",x"f3",x"e7",x"cf",x"99",x"b9",x"ff",
-- [*  *** *]
-- [*  **  *]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [*  **  *]
-- [* ***  *]
-- [********]
x"c3",x"99",x"99",x"c3",x"8b",x"91",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [**    **]
-- [*   * **]
-- [*  *   *]
-- [**     *]
-- [********]
x"e7",x"e7",x"ef",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [*** ****]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"e3",x"cf",x"cf",x"cf",x"cf",x"cf",x"e3",x"ff",
-- [***   **]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [**  ****]
-- [***   **]
-- [********]
x"c7",x"f3",x"f3",x"f3",x"f3",x"f3",x"c7",x"ff",
-- [**   ***]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [****  **]
-- [**   ***]
-- [********]
x"f7",x"d5",x"e3",x"80",x"e3",x"d5",x"f7",x"ff",
-- [**** ***]
-- [** * * *]
-- [***   **]
-- [*       ]
-- [***   **]
-- [** * * *]
-- [**** ***]
-- [********]
x"ff",x"e7",x"e7",x"81",x"e7",x"e7",x"ff",x"ff",
-- [********]
-- [***  ***]
-- [***  ***]
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"e7",x"e7",x"f7",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [***  ***]
-- [***  ***]
-- [**** ***]
-- [********]
x"ff",x"ff",x"ff",x"c3",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [**    **]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"e7",x"e7",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
x"fd",x"f9",x"f3",x"e7",x"cf",x"9f",x"bf",x"ff",
-- [****** *]
-- [*****  *]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [*  *****]
-- [* ******]
-- [********]
x"c3",x"99",x"91",x"81",x"89",x"99",x"c3",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  *   *]
-- [*      *]
-- [*   *  *]
-- [*  **  *]
-- [**    **]
-- [********]
x"e7",x"c7",x"e7",x"e7",x"e7",x"e7",x"81",x"ff",
-- [***  ***]
-- [**   ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [*      *]
-- [********]
x"83",x"99",x"f9",x"e3",x"cf",x"99",x"81",x"ff",
-- [*     **]
-- [*  **  *]
-- [*****  *]
-- [***   **]
-- [**  ****]
-- [*  **  *]
-- [*      *]
-- [********]
x"83",x"99",x"f9",x"f3",x"f9",x"99",x"81",x"ff",
-- [*     **]
-- [*  **  *]
-- [*****  *]
-- [****  **]
-- [*****  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"9f",x"9f",x"93",x"81",x"f3",x"f3",x"f3",x"ff",
-- [*  *****]
-- [*  *****]
-- [*  *  **]
-- [*      *]
-- [****  **]
-- [****  **]
-- [****  **]
-- [********]
x"81",x"99",x"9f",x"83",x"f9",x"99",x"83",x"ff",
-- [*      *]
-- [*  **  *]
-- [*  *****]
-- [*     **]
-- [*****  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"c1",x"99",x"9f",x"83",x"99",x"99",x"c1",x"ff",
-- [**     *]
-- [*  **  *]
-- [*  *****]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"81",x"99",x"f9",x"e1",x"f9",x"f9",x"f9",x"ff",
-- [*      *]
-- [*  **  *]
-- [*****  *]
-- [***    *]
-- [*****  *]
-- [*****  *]
-- [*****  *]
-- [********]
x"c3",x"99",x"99",x"c3",x"99",x"99",x"81",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"c3",x"99",x"99",x"c1",x"f9",x"99",x"83",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [*****  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"ff",x"e7",x"e7",x"ff",x"e7",x"e7",x"ff",x"ff",
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
-- [********]
x"ff",x"e7",x"e7",x"ff",x"e7",x"e7",x"f7",x"ff",
-- [********]
-- [***  ***]
-- [***  ***]
-- [********]
-- [***  ***]
-- [***  ***]
-- [**** ***]
-- [********]
x"ff",x"f3",x"e7",x"cf",x"e7",x"f3",x"ff",x"ff",
-- [********]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [***  ***]
-- [****  **]
-- [********]
-- [********]
x"ff",x"ff",x"c3",x"ff",x"c3",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [**    **]
-- [********]
-- [**    **]
-- [********]
-- [********]
-- [********]
x"ff",x"cf",x"e7",x"f3",x"e7",x"cf",x"ff",x"ff",
-- [********]
-- [**  ****]
-- [***  ***]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [********]
-- [********]
x"81",x"99",x"f9",x"f3",x"e7",x"ff",x"e7",x"ff",
-- [*      *]
-- [*  **  *]
-- [*****  *]
-- [****  **]
-- [***  ***]
-- [********]
-- [***  ***]
-- [********]
x"ff",x"ff",x"ff",x"00",x"00",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
x"c3",x"99",x"99",x"81",x"99",x"99",x"99",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"83",x"99",x"99",x"83",x"99",x"99",x"81",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [********]
x"c3",x"99",x"99",x"9f",x"9f",x"99",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*  *****]
-- [*  *****]
-- [*  **  *]
-- [**     *]
-- [********]
x"83",x"99",x"99",x"99",x"99",x"99",x"83",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"81",x"99",x"9f",x"87",x"9f",x"99",x"81",x"ff",
-- [*      *]
-- [*  **  *]
-- [*  *****]
-- [*    ***]
-- [*  *****]
-- [*  **  *]
-- [*      *]
-- [********]
x"81",x"99",x"9f",x"87",x"9f",x"9f",x"9f",x"ff",
-- [*      *]
-- [*  **  *]
-- [*  *****]
-- [*    ***]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [********]
x"c1",x"99",x"9f",x"91",x"99",x"99",x"c1",x"ff",
-- [**     *]
-- [*  **  *]
-- [*  *****]
-- [*  *   *]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"99",x"99",x"99",x"81",x"99",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"81",x"e7",x"e7",x"e7",x"e7",x"e7",x"81",x"ff",
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [*      *]
-- [********]
x"81",x"99",x"f9",x"f9",x"99",x"99",x"83",x"ff",
-- [*      *]
-- [*  **  *]
-- [*****  *]
-- [*****  *]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [********]
x"99",x"99",x"93",x"87",x"93",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  *  **]
-- [*    ***]
-- [*  *  **]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"9f",x"9f",x"9f",x"9f",x"9f",x"99",x"81",x"ff",
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [*  **  *]
-- [*      *]
-- [********]
x"9c",x"88",x"80",x"80",x"94",x"9c",x"9c",x"ff",
-- [*  ***  ]
-- [*   *   ]
-- [*       ]
-- [*       ]
-- [*  * *  ]
-- [*  ***  ]
-- [*  ***  ]
-- [********]
x"99",x"99",x"89",x"81",x"91",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*   *  *]
-- [*      *]
-- [*  *   *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"c3",x"99",x"99",x"99",x"99",x"99",x"c1",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [**     *]
-- [********]
x"83",x"99",x"99",x"81",x"9f",x"9f",x"9f",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*      *]
-- [*  *****]
-- [*  *****]
-- [*  *****]
-- [********]
x"c3",x"99",x"99",x"99",x"95",x"93",x"c9",x"ff",
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  * * *]
-- [*  *  **]
-- [**  *  *]
-- [********]
x"83",x"99",x"99",x"83",x"99",x"99",x"99",x"ff",
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*     **]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"c1",x"9f",x"8f",x"c3",x"f1",x"f1",x"83",x"ff",
-- [**     *]
-- [*  *****]
-- [*   ****]
-- [**    **]
-- [****   *]
-- [****   *]
-- [*     **]
-- [********]
x"81",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"ff",
-- [*      *]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [********]
x"99",x"99",x"99",x"99",x"99",x"91",x"c3",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [*  *   *]
-- [**    **]
-- [********]
x"99",x"99",x"99",x"d3",x"c3",x"e7",x"e7",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  **  *]
-- [** *  **]
-- [**    **]
-- [***  ***]
-- [***  ***]
-- [********]
x"9c",x"9c",x"94",x"80",x"80",x"88",x"9c",x"ff",
-- [*  ***  ]
-- [*  ***  ]
-- [*  * *  ]
-- [*       ]
-- [*       ]
-- [*   *   ]
-- [*  ***  ]
-- [********]
x"99",x"99",x"c3",x"e7",x"c3",x"99",x"99",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [**    **]
-- [***  ***]
-- [**    **]
-- [*  **  *]
-- [*  **  *]
-- [********]
x"99",x"99",x"91",x"c3",x"e7",x"e7",x"e7",x"ff",
-- [*  **  *]
-- [*  **  *]
-- [*  *   *]
-- [**    **]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [********]
x"81",x"99",x"f3",x"e7",x"cf",x"89",x"81",x"ff",
-- [*      *]
-- [*  **  *]
-- [****  **]
-- [***  ***]
-- [**  ****]
-- [*   *  *]
-- [*      *]
-- [********]
x"e7",x"e7",x"e7",x"00",x"00",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [        ]
-- [        ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"3f",x"3f",x"cf",x"cf",x"3f",x"3f",x"cf",x"cf",
-- [  ******]
-- [  ******]
-- [**  ****]
-- [**  ****]
-- [  ******]
-- [  ******]
-- [**  ****]
-- [**  ****]
x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
x"cc",x"66",x"33",x"99",x"cc",x"66",x"33",x"99",
-- [**  **  ]
-- [ **  ** ]
-- [  **  **]
-- [*  **  *]
-- [**  **  ]
-- [ **  ** ]
-- [  **  **]
-- [*  **  *]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",x"0f",
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
-- [        ]
x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
x"55",x"aa",x"55",x"aa",x"55",x"aa",x"55",x"aa",
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
x"ff",x"ff",x"ff",x"ff",x"55",x"aa",x"55",x"aa",
-- [********]
-- [********]
-- [********]
-- [********]
-- [ * * * *]
-- [* * * * ]
-- [ * * * *]
-- [* * * * ]
x"33",x"66",x"cc",x"99",x"33",x"66",x"cc",x"99",
-- [  **  **]
-- [ **  ** ]
-- [**  **  ]
-- [*  **  *]
-- [  **  **]
-- [ **  ** ]
-- [**  **  ]
-- [*  **  *]
x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
-- [******  ]
x"e7",x"e7",x"e7",x"e0",x"e0",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***     ]
-- [***     ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"ff",x"ff",x"ff",x"ff",x"f0",x"f0",x"f0",x"f0",
-- [********]
-- [********]
-- [********]
-- [********]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
x"e7",x"e7",x"e7",x"e0",x"e0",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [***     ]
-- [***     ]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"07",x"07",x"e7",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [     ***]
-- [     ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
x"ff",x"ff",x"ff",x"e0",x"e0",x"e7",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [***     ]
-- [***     ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"e7",x"e7",x"e7",x"00",x"00",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"00",x"00",x"e7",x"e7",x"e7",
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"e7",x"e7",x"e7",x"07",x"07",x"e7",x"e7",x"e7",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [     ***]
-- [     ***]
-- [***  ***]
-- [***  ***]
-- [***  ***]
x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",x"3f",
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
-- [  ******]
x"1f",x"1f",x"1f",x"1f",x"1f",x"1f",x"1f",x"1f",
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
-- [   *****]
x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
-- [*****   ]
x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"00",x"00",x"00",x"ff",x"ff",x"ff",x"ff",x"ff",
-- [        ]
-- [        ]
-- [        ]
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"ff",x"00",x"00",x"00",
-- [********]
-- [********]
-- [********]
-- [********]
-- [********]
-- [        ]
-- [        ]
-- [        ]
x"ff",x"fe",x"fc",x"b9",x"93",x"c7",x"ef",x"ff",
-- [********]
-- [******* ]
-- [******  ]
-- [* ***  *]
-- [*  *  **]
-- [**   ***]
-- [*** ****]
-- [********]
x"ff",x"ff",x"ff",x"ff",x"0f",x"0f",x"0f",x"0f",
-- [********]
-- [********]
-- [********]
-- [********]
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
x"f0",x"f0",x"f0",x"f0",x"ff",x"ff",x"ff",x"ff",
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
-- [********]
-- [********]
-- [********]
-- [********]
x"e7",x"e7",x"e7",x"07",x"07",x"ff",x"ff",x"ff",
-- [***  ***]
-- [***  ***]
-- [***  ***]
-- [     ***]
-- [     ***]
-- [********]
-- [********]
-- [********]
x"0f",x"0f",x"0f",x"0f",x"ff",x"ff",x"ff",x"ff",
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [********]
-- [********]
-- [********]
-- [********]
x"0f",x"0f",x"0f",x"0f",x"f0",x"f0",x"f0",x"f0" 
-- [    ****]
-- [    ****]
-- [    ****]
-- [    ****]
-- [****    ]
-- [****    ]
-- [****    ]
-- [****    ]
);

begin

--process for read and write operation.
PROCESS(Clk,ram,writeclk)
BEGIN

  if(rising_edge(writeClk)) then 
    if writecs='1' then
      if(we='1') then
        ram(to_integer(writeaddress)) <= data_i;
      end if;
    end if;
    data_o <= ram(address);
  end if;
END PROCESS;

end Behavioral;
