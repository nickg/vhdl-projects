library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

--
entity hyppo is
  port (Clk : in std_logic;
        address : in std_logic_vector(13 downto 0);
        address_i : in std_logic_vector(13 downto 0);
        -- Yes, we do have a write enable, because we allow modification of ROMs
        -- in the running machine, unless purposely disabled.  This gives us
        -- something like the WOM that the Amiga had.
        we : in std_logic;
        -- chip select, active low       
        cs : in std_logic;
        data_i : in std_logic_vector(7 downto 0);
        data_o : out std_logic_vector(7 downto 0)
        );
end hyppo;

architecture Behavioral of hyppo is

-- 16K x 8bit pre-initialised RAM
  type ram_t is array (0 to 16383) of std_logic_vector(7 downto 0);
  signal ram : ram_t := (x"4C",x"B9",x"8B",x"EA",x"4C",x"AD",x"9D",x"EA",x"4C",x"08",x"86",x"EA",x"4C",x"FC",x"AD",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"CF",x"9F",x"EA",x"4C",x"DC",x"9F",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"BB",x"9F",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"1F",x"9F",x"EA",x"4C",x"BA",x"A3",x"EA",x"4C",x"55",x"9D",x"EA",x"4C",x"1F",x"9F",x"EA",x"4C",x"C4",x"9F",x"EA",x"4C",x"26",x"A1",x"EA",x"4C",x"69",x"A1",x"EA",x"4C",x"1F",x"9F",x"EA",x"4C",x"1F",x"9F",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"4C",x"00",x"82",x"EA",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BA",x"A3",x"A4",x"AB",x"BA",x"A3",x"A4",x"AB",x"AD",x"47",x"D6",x"29",x"FE",x"8D",x"47",x"D6",x"A9",x"FF",x"8D",x"40",x"D6",x"8D",x"7F",x"D6",x"AD",x"F8",x"BC",x"8D",x"40",x"D6",x"20",x"CA",x"A0",x"AD",x"47",x"D6",x"09",x"01",x"8D",x"47",x"D6",x"8D",x"7F",x"D6",x"20",x"CA",x"A0",x"8D",x"40",x"D6",x"AD",x"47",x"D6",x"29",x"FE",x"8D",x"47",x"D6",x"8D",x"7F",x"D6",x"4C",x"00",x"82",x"0A",x"80",x"00",x"81",x"00",x"00",x"00",x"FF",x"77",x"00",x"00",x"04",x"FF",x"07",x"00",x"00",x"00",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"82",x"8D",x"01",x"D7",x"A9",x"38",x"8D",x"05",x"D7",x"4C",x"C5",x"AC",x"A2",x"03",x"BD",x"C0",x"BB",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"A9",x"01",x"8D",x"FC",x"BC",x"20",x"D3",x"A0",x"90",x"7F",x"A9",x"42",x"8D",x"FC",x"BC",x"A2",x"0A",x"BD",x"00",x"DE",x"DD",x"7D",x"85",x"D0",x"70",x"CA",x"10",x"F5",x"A9",x"00",x"8D",x"FC",x"BC",x"A2",x"10",x"BD",x"00",x"DE",x"9D",x"C0",x"BB",x"E8",x"E0",x"30",x"D0",x"F5",x"A2",x"C0",x"A0",x"85",x"20",x"2B",x"A9",x"A0",x"00",x"AB",x"DD",x"BB",x"20",x"A4",x"A9",x"AB",x"DC",x"BB",x"20",x"A4",x"A9",x"AB",x"ED",x"BB",x"20",x"A4",x"A9",x"AB",x"EC",x"BB",x"20",x"A4",x"A9",x"AB",x"DB",x"BB",x"20",x"A4",x"A9",x"AB",x"DA",x"BB",x"20",x"A4",x"A9",x"AB",x"D9",x"BB",x"20",x"A4",x"A9",x"AB",x"D8",x"BB",x"20",x"A4",x"A9",x"A9",x"01",x"8D",x"FD",x"BC",x"A2",x"AC",x"A0",x"85",x"20",x"2B",x"A9",x"20",x"04",x"84",x"AD",x"0E",x"DE",x"10",x"21",x"20",x"14",x"84",x"B0",x"07",x"A2",x"E4",x"A0",x"85",x"20",x"2B",x"A9",x"38",x"60",x"A2",x"88",x"A0",x"85",x"20",x"2B",x"A9",x"A0",x"00",x"AB",x"FC",x"BC",x"20",x"A4",x"A9",x"A3",x"00",x"18",x"60",x"AD",x"07",x"A4",x"C9",x"4C",x"F0",x"D8",x"4C",x"49",x"82",x"20",x"04",x"84",x"8D",x"7F",x"D6",x"20",x"0A",x"84",x"8D",x"7F",x"D6",x"20",x"F7",x"83",x"8D",x"7F",x"D6",x"20",x"14",x"84",x"8D",x"7F",x"D6",x"AE",x"41",x"D6",x"20",x"64",x"83",x"20",x"B1",x"86",x"AD",x"00",x"BD",x"C9",x"FF",x"D0",x"05",x"A9",x"00",x"8D",x"00",x"BD",x"A9",x"FF",x"CD",x"12",x"D0",x"D0",x"FB",x"CE",x"19",x"D0",x"8D",x"7F",x"D6",x"AE",x"DC",x"BB",x"8E",x"41",x"D6",x"AC",x"DD",x"BB",x"8C",x"42",x"D6",x"4C",x"16",x"82",x"AE",x"41",x"D6",x"AC",x"42",x"D6",x"20",x"64",x"83",x"8D",x"7F",x"D6",x"DA",x"5A",x"AD",x"FD",x"BC",x"D0",x"07",x"A9",x"FF",x"8D",x"FC",x"BC",x"18",x"60",x"CC",x"DD",x"BB",x"F0",x"02",x"90",x"0E",x"EC",x"DC",x"BB",x"F0",x"02",x"90",x"07",x"A9",x"02",x"8D",x"FC",x"BC",x"18",x"60",x"20",x"B9",x"83",x"A2",x"03",x"BD",x"D8",x"BB",x"9D",x"70",x"D7",x"CA",x"10",x"F7",x"FA",x"8E",x"74",x"D7",x"7A",x"8C",x"75",x"D7",x"A9",x"00",x"8D",x"76",x"D7",x"8D",x"77",x"D7",x"A2",x"00",x"A0",x"03",x"18",x"BD",x"78",x"D7",x"7D",x"81",x"D6",x"9D",x"81",x"D6",x"E8",x"88",x"10",x"F3",x"38",x"60",x"AD",x"C0",x"BB",x"18",x"6D",x"D0",x"BB",x"8D",x"81",x"D6",x"A2",x"01",x"BD",x"C0",x"BB",x"7D",x"D0",x"BB",x"9D",x"81",x"D6",x"E8",x"E0",x"04",x"D0",x"F2",x"AD",x"81",x"D6",x"18",x"6D",x"DE",x"BB",x"8D",x"81",x"D6",x"AD",x"82",x"D6",x"6D",x"DF",x"BB",x"8D",x"82",x"D6",x"AD",x"83",x"D6",x"69",x"00",x"8D",x"83",x"D6",x"AD",x"84",x"D6",x"69",x"00",x"8D",x"84",x"D6",x"60",x"A2",x"03",x"A9",x"00",x"9D",x"81",x"D6",x"CA",x"10",x"FA",x"4C",x"13",x"A1",x"20",x"F7",x"83",x"4C",x"D3",x"A0",x"20",x"F7",x"83",x"20",x"44",x"A0",x"38",x"60",x"18",x"60",x"AD",x"00",x"DE",x"C9",x"01",x"D0",x"F7",x"AD",x"01",x"DE",x"C9",x"01",x"D0",x"F0",x"AD",x"20",x"DE",x"8D",x"03",x"D7",x"A9",x"28",x"1C",x"54",x"D0",x"2D",x"21",x"DE",x"0C",x"54",x"D0",x"AE",x"58",x"D0",x"AD",x"6F",x"D0",x"29",x"3F",x"8D",x"6F",x"D0",x"AD",x"02",x"DE",x"29",x"C0",x"0D",x"6F",x"D0",x"8D",x"6F",x"D0",x"8D",x"E4",x"A7",x"8E",x"58",x"D0",x"AD",x"02",x"DE",x"29",x"80",x"D0",x"12",x"AD",x"0E",x"DC",x"09",x"80",x"8D",x"0E",x"DC",x"AD",x"0E",x"DD",x"09",x"80",x"8D",x"0E",x"DD",x"80",x"10",x"AD",x"0E",x"DC",x"29",x"7F",x"8D",x"0E",x"DC",x"AD",x"0E",x"DD",x"29",x"7F",x"8D",x"0E",x"DD",x"AD",x"0D",x"DE",x"8D",x"1A",x"D6",x"A9",x"00",x"8D",x"3C",x"D6",x"AD",x"22",x"DE",x"F0",x"05",x"A9",x"0F",x"8D",x"3C",x"D6",x"AD",x"0C",x"DE",x"A3",x"00",x"A9",x"07",x"8D",x"13",x"BF",x"A2",x"FE",x"8E",x"12",x"BF",x"E8",x"8E",x"11",x"BF",x"8E",x"10",x"BF",x"EA",x"92",x"10",x"AD",x"03",x"DE",x"29",x"01",x"8D",x"FE",x"D6",x"AD",x"03",x"DE",x"29",x"40",x"F0",x"06",x"20",x"DA",x"A1",x"4C",x"CB",x"84",x"AD",x"03",x"DE",x"29",x"20",x"D0",x"06",x"20",x"55",x"A2",x"4C",x"CB",x"84",x"20",x"5F",x"A2",x"AD",x"04",x"DE",x"8D",x"A1",x"D6",x"AD",x"05",x"DE",x"8D",x"1B",x"D6",x"A9",x"4C",x"8D",x"D1",x"94",x"AD",x"0F",x"DE",x"10",x"05",x"A9",x"2C",x"8D",x"D1",x"94",x"A2",x"05",x"BD",x"06",x"DE",x"9D",x"E9",x"D6",x"CA",x"10",x"F7",x"AD",x"10",x"DE",x"F0",x"0B",x"A2",x"0F",x"BD",x"10",x"DE",x"9D",x"1C",x"B3",x"CA",x"10",x"F7",x"38",x"60",x"20",x"09",x"85",x"8D",x"7F",x"D6",x"A9",x"16",x"8D",x"10",x"BF",x"A9",x"00",x"8D",x"11",x"BF",x"8D",x"13",x"BF",x"A9",x"02",x"8D",x"12",x"BF",x"A3",x"00",x"EA",x"B2",x"10",x"C9",x"56",x"F0",x"01",x"60",x"1B",x"EA",x"B2",x"10",x"C9",x"39",x"D0",x"34",x"1B",x"EA",x"B2",x"10",x"C9",x"30",x"F0",x"3A",x"C9",x"31",x"D0",x"28",x"1B",x"EA",x"B2",x"10",x"C9",x"30",x"D0",x"20",x"1B",x"EA",x"B2",x"10",x"C9",x"36",x"B0",x"18",x"C9",x"35",x"90",x"22",x"1B",x"EA",x"B2",x"10",x"C9",x"32",x"90",x"1A",x"C9",x"33",x"B0",x"08",x"1B",x"EA",x"B2",x"10",x"C9",x"33",x"90",x"0E",x"A3",x"00",x"A9",x"01",x"0C",x"03",x"D7",x"A2",x"C4",x"A0",x"B2",x"4C",x"2B",x"A9",x"A3",x"00",x"A9",x"01",x"1C",x"03",x"D7",x"A2",x"B2",x"A0",x"B2",x"4C",x"2B",x"A9",x"4D",x"45",x"47",x"41",x"36",x"35",x"53",x"59",x"53",x"30",x"30",x"53",x"59",x"53",x"54",x"45",x"4D",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"45",x"52",x"52",x"4F",x"52",x"3A",x"20",x"28",x"45",x"52",x"52",x"4E",x"4F",x"3A",x"20",x"24",x"24",x"29",x"00",x"53",x"59",x"53",x"54",x"45",x"4D",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"4F",x"4B",x"00",x"53",x"59",x"53",x"3A",x"20",x"24",x"24",x"24",x"24",x"20",x"46",x"52",x"5A",x"20",x"2B",x"20",x"24",x"24",x"24",x"24",x"20",x"53",x"56",x"43",x"20",x"58",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"53",x"59",x"53",x"50",x"41",x"52",x"54",x"20",x"43",x"4F",x"4E",x"46",x"49",x"47",x"20",x"49",x"4E",x"56",x"41",x"4C",x"49",x"44",x"2E",x"20",x"50",x"4C",x"45",x"41",x"53",x"45",x"20",x"53",x"45",x"54",x"2E",x"00",x"78",x"D8",x"29",x"FE",x"AA",x"7C",x"10",x"86",x"0F",x"83",x"15",x"83",x"21",x"83",x"1B",x"83",x"03",x"85",x"35",x"82",x"35",x"82",x"35",x"82",x"58",x"83",x"27",x"83",x"01",x"8B",x"49",x"83",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"20",x"64",x"83",x"B0",x"01",x"60",x"20",x"93",x"8A",x"20",x"4E",x"87",x"A2",x"00",x"20",x"BB",x"87",x"8A",x"18",x"69",x"08",x"AA",x"BD",x"24",x"8B",x"C9",x"FF",x"D0",x"F1",x"20",x"AA",x"87",x"60",x"20",x"13",x"A1",x"A2",x"00",x"20",x"5E",x"A0",x"20",x"B1",x"88",x"A9",x"47",x"8D",x"2F",x"D0",x"A9",x"53",x"8D",x"2F",x"D0",x"8A",x"18",x"69",x"08",x"AA",x"BD",x"24",x"8B",x"C9",x"FF",x"D0",x"E4",x"20",x"BC",x"99",x"AE",x"13",x"BD",x"F0",x"27",x"A2",x"00",x"BD",x"15",x"BD",x"9D",x"67",x"BC",x"E8",x"EC",x"13",x"BD",x"D0",x"F4",x"A9",x"00",x"9D",x"67",x"BC",x"8E",x"66",x"BC",x"AD",x"11",x"BD",x"29",x"04",x"48",x"20",x"CE",x"99",x"68",x"C9",x"00",x"F0",x"03",x"20",x"E6",x"8F",x"AE",x"14",x"BD",x"F0",x"27",x"A2",x"00",x"BD",x"35",x"BD",x"9D",x"67",x"BC",x"E8",x"EC",x"14",x"BD",x"D0",x"F4",x"A9",x"00",x"9D",x"67",x"BC",x"8E",x"66",x"BC",x"AD",x"12",x"BD",x"29",x"04",x"48",x"20",x"4F",x"9A",x"68",x"C9",x"00",x"F0",x"03",x"20",x"E6",x"8F",x"A9",x"0F",x"8D",x"18",x"D4",x"8D",x"38",x"D4",x"8D",x"58",x"D4",x"8D",x"78",x"D4",x"60",x"20",x"5E",x"A0",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"55",x"A0",x"90",x"F3",x"20",x"13",x"A1",x"38",x"60",x"EE",x"20",x"D0",x"A9",x"00",x"8D",x"B9",x"87",x"8D",x"BA",x"87",x"20",x"5E",x"A0",x"20",x"3E",x"A0",x"A9",x"04",x"8D",x"80",x"D6",x"20",x"55",x"A0",x"4C",x"74",x"87",x"EE",x"B9",x"87",x"D0",x"EA",x"EE",x"BA",x"87",x"D0",x"E5",x"CE",x"20",x"D0",x"20",x"13",x"A1",x"38",x"60",x"EE",x"20",x"D0",x"A9",x"00",x"8D",x"B9",x"87",x"8D",x"BA",x"87",x"20",x"5E",x"A0",x"20",x"3E",x"A0",x"A9",x"05",x"8D",x"80",x"D6",x"20",x"55",x"A0",x"4C",x"A2",x"87",x"EE",x"B9",x"87",x"D0",x"EA",x"EE",x"BA",x"87",x"D0",x"E5",x"CE",x"20",x"D0",x"20",x"13",x"A1",x"38",x"60",x"20",x"55",x"A0",x"20",x"3E",x"A0",x"A9",x"06",x"8D",x"80",x"D6",x"20",x"55",x"A0",x"60",x"00",x"00",x"BD",x"24",x"8B",x"C9",x"FF",x"D0",x"01",x"60",x"DA",x"AA",x"20",x"71",x"89",x"FA",x"BD",x"1D",x"8B",x"8D",x"C6",x"8A",x"BD",x"1E",x"8B",x"8D",x"C7",x"8A",x"BD",x"1F",x"8B",x"4A",x"4A",x"4A",x"4A",x"8D",x"BF",x"8A",x"BD",x"20",x"8B",x"0A",x"0A",x"0A",x"0A",x"0D",x"BF",x"8A",x"8D",x"BF",x"8A",x"BD",x"1F",x"8B",x"29",x"0F",x"8D",x"C8",x"8A",x"A9",x"00",x"8D",x"C9",x"8A",x"A9",x"6E",x"8D",x"CA",x"8A",x"A9",x"0D",x"8D",x"CB",x"8A",x"A9",x"FF",x"8D",x"C1",x"8A",x"BD",x"21",x"8B",x"8D",x"B5",x"8B",x"BD",x"22",x"8B",x"8D",x"B6",x"8B",x"BD",x"23",x"8B",x"29",x"7F",x"8D",x"B7",x"8B",x"20",x"8F",x"88",x"0D",x"B5",x"8B",x"0D",x"B7",x"8B",x"F0",x"3C",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"8A",x"8D",x"01",x"D7",x"A9",x"BD",x"8D",x"05",x"D7",x"EE",x"20",x"D0",x"20",x"7C",x"87",x"CE",x"20",x"D0",x"20",x"64",x"88",x"F0",x"1C",x"20",x"73",x"88",x"20",x"64",x"88",x"F0",x"14",x"AD",x"C7",x"8A",x"18",x"69",x"02",x"8D",x"C7",x"8A",x"AD",x"C8",x"8A",x"69",x"00",x"8D",x"C8",x"8A",x"4C",x"1C",x"88",x"60",x"AD",x"B7",x"8B",x"30",x"07",x"0D",x"B6",x"8B",x"0D",x"B5",x"8B",x"60",x"A9",x"00",x"60",x"38",x"AD",x"B5",x"8B",x"ED",x"C4",x"8A",x"8D",x"B5",x"8B",x"AD",x"B6",x"8B",x"ED",x"C5",x"8A",x"8D",x"B6",x"8B",x"AD",x"B7",x"8B",x"E9",x"00",x"8D",x"B7",x"8B",x"60",x"AD",x"B6",x"8B",x"29",x"FE",x"0D",x"B7",x"8B",x"F0",x"0B",x"A9",x"00",x"8D",x"C4",x"8A",x"A9",x"02",x"8D",x"C5",x"8A",x"60",x"AD",x"B5",x"8B",x"8D",x"C4",x"8A",x"AD",x"B6",x"8B",x"8D",x"C5",x"8A",x"60",x"BD",x"24",x"8B",x"C9",x"FF",x"F0",x"04",x"C5",x"0C",x"D0",x"01",x"60",x"DA",x"AA",x"20",x"74",x"89",x"FA",x"BD",x"1D",x"8B",x"8D",x"C9",x"8A",x"BD",x"1E",x"8B",x"8D",x"CA",x"8A",x"BD",x"1F",x"8B",x"4A",x"4A",x"4A",x"4A",x"8D",x"C1",x"8A",x"BD",x"20",x"8B",x"0A",x"0A",x"0A",x"0A",x"0D",x"C1",x"8A",x"8D",x"C1",x"8A",x"BD",x"1F",x"8B",x"29",x"0F",x"8D",x"CB",x"8A",x"A9",x"00",x"8D",x"C6",x"8A",x"A9",x"6E",x"8D",x"C7",x"8A",x"A9",x"0D",x"8D",x"C8",x"8A",x"A9",x"FF",x"8D",x"BF",x"8A",x"BD",x"21",x"8B",x"8D",x"B5",x"8B",x"BD",x"22",x"8B",x"8D",x"B6",x"8B",x"BD",x"23",x"8B",x"8D",x"B8",x"8B",x"29",x"7F",x"8D",x"B7",x"8B",x"EE",x"20",x"D0",x"20",x"3C",x"87",x"CE",x"20",x"D0",x"20",x"8F",x"88",x"0D",x"B5",x"8B",x"0D",x"B7",x"8B",x"F0",x"38",x"2C",x"B8",x"8B",x"30",x"12",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"8A",x"8D",x"01",x"D7",x"A9",x"BD",x"8D",x"05",x"D7",x"20",x"64",x"88",x"F0",x"1C",x"20",x"73",x"88",x"20",x"64",x"88",x"F0",x"14",x"AD",x"CA",x"8A",x"18",x"69",x"02",x"8D",x"CA",x"8A",x"AD",x"CB",x"8A",x"69",x"00",x"8D",x"CB",x"8A",x"4C",x"19",x"89",x"DA",x"48",x"BD",x"24",x"8B",x"AA",x"20",x"77",x"89",x"68",x"FA",x"60",x"7C",x"44",x"8A",x"7C",x"54",x"8A",x"7C",x"66",x"8A",x"A9",x"00",x"85",x"00",x"A9",x"62",x"85",x"01",x"A9",x"FD",x"85",x"02",x"A9",x"0F",x"85",x"03",x"A3",x"8F",x"6B",x"AA",x"EA",x"B2",x"00",x"E0",x"00",x"F0",x"0B",x"E0",x"80",x"F0",x"07",x"E0",x"85",x"F0",x"03",x"9D",x"80",x"D6",x"CA",x"3B",x"C2",x"FF",x"D0",x"E6",x"A3",x"00",x"60",x"A9",x"00",x"85",x"00",x"A9",x"10",x"85",x"01",x"A0",x"00",x"A2",x"10",x"A9",x"40",x"8D",x"10",x"BF",x"A9",x"26",x"8D",x"11",x"BF",x"A9",x"FD",x"8D",x"12",x"BF",x"A9",x"0F",x"8D",x"13",x"BF",x"A3",x"00",x"EA",x"B2",x"10",x"A9",x"41",x"8D",x"10",x"BF",x"EA",x"B2",x"10",x"91",x"00",x"C8",x"D0",x"F8",x"E6",x"01",x"CA",x"D0",x"F3",x"60",x"A9",x"00",x"85",x"00",x"A9",x"62",x"85",x"01",x"A9",x"FD",x"85",x"02",x"A9",x"0F",x"85",x"03",x"A3",x"8F",x"6B",x"AA",x"BD",x"80",x"D6",x"EA",x"92",x"00",x"CA",x"3B",x"C2",x"FF",x"D0",x"F2",x"A3",x"00",x"A9",x"FF",x"8D",x"BF",x"8A",x"8D",x"C1",x"8A",x"A9",x"8D",x"8D",x"C8",x"8A",x"8D",x"CB",x"8A",x"A9",x"00",x"8D",x"C6",x"8A",x"A9",x"6E",x"8D",x"C7",x"8A",x"A9",x"00",x"8D",x"C9",x"8A",x"A9",x"60",x"8D",x"CA",x"8A",x"A9",x"00",x"8D",x"C4",x"8A",x"A9",x"02",x"8D",x"C5",x"8A",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"8A",x"8D",x"01",x"D7",x"A9",x"BD",x"8D",x"05",x"D7",x"60",x"43",x"8A",x"CE",x"8A",x"CE",x"8A",x"CE",x"8A",x"CE",x"8A",x"E1",x"89",x"A9",x"89",x"B6",x"8A",x"78",x"8A",x"CE",x"8A",x"CE",x"8A",x"CE",x"8A",x"CE",x"8A",x"78",x"8A",x"78",x"8A",x"78",x"8A",x"78",x"8A",x"79",x"8A",x"78",x"8A",x"78",x"8A",x"78",x"8A",x"78",x"8A",x"78",x"8A",x"78",x"8A",x"78",x"8A",x"7A",x"8A",x"60",x"60",x"A9",x"11",x"85",x"00",x"A9",x"6E",x"85",x"01",x"A9",x"FD",x"85",x"02",x"A9",x"0F",x"85",x"03",x"A3",x"00",x"EA",x"B2",x"00",x"8D",x"51",x"D6",x"60",x"A2",x"0F",x"BD",x"80",x"D6",x"9D",x"A5",x"8A",x"CA",x"10",x"F7",x"AD",x"70",x"D0",x"8D",x"B5",x"8A",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"B5",x"8A",x"8D",x"70",x"D0",x"60",x"0A",x"80",x"00",x"81",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"8A",x"18",x"E9",x"02",x"0A",x"0A",x"0A",x"0A",x"0A",x"09",x"3F",x"8D",x"70",x"D0",x"60",x"AD",x"11",x"D6",x"F0",x"FB",x"AD",x"11",x"D6",x"D0",x"FB",x"60",x"AD",x"81",x"D6",x"8D",x"00",x"08",x"AD",x"82",x"D6",x"8D",x"01",x"08",x"AD",x"83",x"D6",x"8D",x"02",x"08",x"AD",x"84",x"D6",x"8D",x"03",x"08",x"60",x"AE",x"41",x"D6",x"86",x"00",x"AD",x"42",x"D6",x"29",x"7F",x"85",x"01",x"A2",x"98",x"A0",x"00",x"B9",x"1D",x"8B",x"91",x"00",x"C8",x"CA",x"D0",x"F7",x"4C",x"16",x"82",x"A5",x"8A",x"FF",x"0F",x"10",x"00",x"00",x"00",x"00",x"60",x"FD",x"0F",x"90",x"00",x"00",x"0A",x"00",x"6C",x"FD",x"0F",x"00",x"02",x"00",x"00",x"00",x"BD",x"FF",x"0F",x"00",x"01",x"00",x"00",x"40",x"36",x"FD",x"0F",x"3E",x"00",x"00",x"10",x"00",x"31",x"FD",x"0F",x"00",x"03",x"00",x"02",x"00",x"31",x"FD",x"0F",x"00",x"03",x"00",x"04",x"00",x"31",x"FD",x"0F",x"00",x"03",x"00",x"06",x"00",x"31",x"FD",x"0F",x"00",x"03",x"00",x"08",x"00",x"00",x"F8",x"0F",x"00",x"80",x"00",x"00",x"00",x"3C",x"FD",x"0F",x"00",x"02",x"00",x"00",x"00",x"30",x"FD",x"0F",x"80",x"00",x"00",x"0E",x"30",x"00",x"FD",x"0F",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"BD",x"00",x"00",x"00",x"01",x"00",x"00",x"10",x"37",x"FD",x"0F",x"F0",x"00",x"00",x"00",x"00",x"B0",x"FD",x"0F",x"00",x"50",x"00",x"00",x"00",x"10",x"00",x"00",x"00",x"10",x"80",x"0C",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"78",x"D8",x"29",x"7E",x"AA",x"7C",x"C1",x"8B",x"86",x"8C",x"9D",x"8C",x"FB",x"8C",x"A6",x"8C",x"02",x"90",x"02",x"90",x"63",x"8F",x"02",x"90",x"02",x"90",x"15",x"8F",x"23",x"8F",x"51",x"8F",x"71",x"8F",x"54",x"8F",x"02",x"90",x"04",x"8D",x"7F",x"8F",x"B4",x"8C",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"DC",x"8C",x"A1",x"8F",x"AC",x"8F",x"9B",x"8F",x"BD",x"8C",x"B2",x"8F",x"D6",x"8C",x"5A",x"8F",x"BA",x"8C",x"BB",x"8F",x"C7",x"8F",x"CD",x"8F",x"C1",x"8F",x"D3",x"8F",x"35",x"82",x"35",x"82",x"35",x"82",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"35",x"82",x"35",x"82",x"35",x"82",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"02",x"90",x"78",x"8C",x"6D",x"8C",x"47",x"8C",x"5A",x"8C",x"35",x"82",x"35",x"82",x"41",x"8C",x"BA",x"A3",x"8C",x"7C",x"D6",x"4C",x"16",x"82",x"20",x"A6",x"AB",x"90",x"0B",x"A0",x"05",x"B9",x"4A",x"D6",x"91",x"06",x"88",x"10",x"F8",x"38",x"4C",x"AC",x"8C",x"20",x"A6",x"AB",x"90",x"0B",x"A0",x"05",x"B1",x"06",x"99",x"4A",x"D6",x"88",x"10",x"F8",x"38",x"4C",x"AC",x"8C",x"AD",x"7D",x"D6",x"49",x"20",x"8D",x"7D",x"D6",x"4C",x"80",x"8C",x"AD",x"7D",x"D6",x"49",x"04",x"8D",x"7D",x"D6",x"8D",x"40",x"D6",x"4C",x"16",x"82",x"A9",x"02",x"8D",x"41",x"D6",x"A9",x"01",x"8D",x"40",x"D6",x"A9",x"01",x"8D",x"42",x"D6",x"A9",x"02",x"8D",x"43",x"D6",x"4C",x"16",x"82",x"AD",x"02",x"BC",x"8D",x"40",x"D6",x"4C",x"16",x"82",x"AE",x"41",x"D6",x"20",x"B6",x"92",x"B0",x"03",x"4C",x"24",x"82",x"4C",x"16",x"82",x"20",x"05",x"90",x"4C",x"16",x"82",x"A9",x"08",x"2C",x"A9",x"00",x"85",x"1B",x"AD",x"41",x"D6",x"85",x"18",x"AD",x"42",x"D6",x"85",x"19",x"AD",x"43",x"D6",x"85",x"1A",x"20",x"99",x"98",x"4C",x"AC",x"8C",x"20",x"A6",x"AB",x"4C",x"AC",x"8C",x"20",x"A6",x"AB",x"90",x"0C",x"A6",x"06",x"A4",x"07",x"20",x"9C",x"99",x"90",x"03",x"4C",x"16",x"82",x"8D",x"FB",x"BC",x"4C",x"24",x"82",x"A9",x"11",x"8D",x"FB",x"BC",x"4C",x"24",x"82",x"AD",x"03",x"BC",x"8D",x"40",x"D6",x"4C",x"16",x"82",x"20",x"DE",x"93",x"90",x"09",x"18",x"A9",x"8D",x"8D",x"FB",x"BC",x"4C",x"24",x"82",x"AD",x"43",x"D6",x"4A",x"4A",x"4A",x"18",x"69",x"01",x"8D",x"04",x"BF",x"A9",x"80",x"85",x"10",x"A9",x"00",x"85",x"11",x"85",x"12",x"85",x"13",x"A9",x"00",x"8D",x"05",x"BF",x"20",x"BE",x"A0",x"A2",x"03",x"B5",x"10",x"9D",x"B3",x"BC",x"CA",x"10",x"F8",x"20",x"04",x"8F",x"A2",x"00",x"BD",x"00",x"DE",x"D0",x"08",x"BD",x"00",x"DF",x"D0",x"03",x"E8",x"D0",x"F3",x"F0",x"08",x"A9",x"00",x"8D",x"05",x"BF",x"4C",x"63",x"8D",x"EE",x"05",x"BF",x"AD",x"05",x"BF",x"CD",x"04",x"BF",x"F0",x"1C",x"A9",x"80",x"18",x"65",x"10",x"85",x"10",x"A5",x"11",x"69",x"00",x"85",x"11",x"A5",x"12",x"69",x"00",x"85",x"12",x"A5",x"13",x"69",x"00",x"85",x"13",x"4C",x"32",x"8D",x"CE",x"05",x"BF",x"AD",x"05",x"BF",x"F0",x"1F",x"A5",x"10",x"38",x"E9",x"80",x"85",x"10",x"A5",x"11",x"E9",x"00",x"85",x"11",x"A5",x"12",x"E9",x"00",x"85",x"12",x"A5",x"13",x"E9",x"00",x"85",x"13",x"CE",x"05",x"BF",x"4C",x"82",x"8D",x"20",x"C1",x"8E",x"B0",x"01",x"60",x"A0",x"1F",x"A9",x"00",x"91",x"00",x"C0",x"0B",x"D0",x"02",x"A9",x"20",x"88",x"10",x"F5",x"A0",x"00",x"A2",x"00",x"BD",x"67",x"BC",x"C9",x"2E",x"D0",x"04",x"A0",x"07",x"D0",x"06",x"C9",x"00",x"F0",x"0A",x"91",x"00",x"F0",x"06",x"E8",x"C8",x"C0",x"0B",x"D0",x"E7",x"A0",x"0B",x"A9",x"20",x"91",x"00",x"A0",x"1A",x"A5",x"10",x"91",x"00",x"C8",x"A5",x"11",x"91",x"00",x"A0",x"14",x"A5",x"12",x"91",x"00",x"C8",x"A5",x"13",x"91",x"00",x"A0",x"1C",x"AD",x"41",x"D6",x"91",x"00",x"C8",x"AD",x"42",x"D6",x"91",x"00",x"C8",x"AD",x"43",x"D6",x"91",x"00",x"C8",x"A9",x"00",x"91",x"00",x"20",x"44",x"A0",x"20",x"55",x"A0",x"AD",x"04",x"BF",x"8D",x"05",x"BF",x"A2",x"03",x"B5",x"10",x"9D",x"B3",x"BC",x"CA",x"10",x"F8",x"20",x"04",x"8F",x"A0",x"00",x"A5",x"10",x"18",x"69",x"01",x"85",x"10",x"99",x"00",x"DE",x"C8",x"A5",x"11",x"69",x"00",x"85",x"11",x"99",x"00",x"DE",x"C8",x"A5",x"12",x"69",x"00",x"85",x"12",x"99",x"00",x"DE",x"C8",x"A5",x"13",x"69",x"00",x"85",x"13",x"99",x"00",x"DE",x"C8",x"D0",x"D5",x"A5",x"10",x"18",x"69",x"01",x"85",x"10",x"99",x"00",x"DF",x"C8",x"A5",x"11",x"69",x"00",x"85",x"11",x"99",x"00",x"DF",x"C8",x"A5",x"12",x"69",x"00",x"85",x"12",x"99",x"00",x"DF",x"C8",x"A5",x"13",x"69",x"00",x"85",x"13",x"99",x"00",x"DF",x"C8",x"D0",x"D5",x"AD",x"05",x"BF",x"C9",x"01",x"D0",x"12",x"A9",x"F8",x"8D",x"FC",x"DF",x"A9",x"FF",x"8D",x"FD",x"DF",x"8D",x"FE",x"DF",x"A9",x"0F",x"8D",x"FF",x"DF",x"20",x"44",x"A0",x"20",x"55",x"A0",x"AD",x"04",x"BC",x"09",x"09",x"A8",x"A2",x"00",x"BD",x"81",x"D6",x"79",x"00",x"BB",x"C8",x"E8",x"E0",x"04",x"D0",x"F4",x"20",x"44",x"A0",x"20",x"55",x"A0",x"CE",x"05",x"BF",x"F0",x"03",x"4C",x"18",x"8E",x"4C",x"16",x"82",x"20",x"0A",x"94",x"20",x"BE",x"A0",x"20",x"34",x"97",x"A2",x"00",x"A9",x"DE",x"85",x"01",x"BD",x"00",x"DE",x"C9",x"00",x"F0",x"29",x"C9",x"E5",x"F0",x"25",x"8A",x"69",x"20",x"AA",x"D0",x"EF",x"E6",x"01",x"BD",x"00",x"DE",x"C9",x"00",x"F0",x"16",x"C9",x"E5",x"F0",x"12",x"8A",x"69",x"20",x"AA",x"D0",x"EF",x"20",x"51",x"97",x"B0",x"CE",x"A9",x"8E",x"8D",x"FB",x"BC",x"18",x"60",x"86",x"00",x"38",x"60",x"20",x"54",x"98",x"A2",x"03",x"BD",x"B3",x"BC",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"4C",x"D3",x"A0",x"20",x"0A",x"94",x"B0",x"06",x"AD",x"FB",x"BC",x"4C",x"24",x"82",x"4C",x"10",x"82",x"20",x"BE",x"A0",x"AE",x"41",x"D6",x"8E",x"F8",x"BC",x"20",x"0D",x"97",x"90",x"1A",x"8D",x"F9",x"BC",x"20",x"45",x"94",x"90",x"12",x"20",x"A6",x"AB",x"90",x"0D",x"A0",x"56",x"B9",x"0F",x"BC",x"91",x"06",x"88",x"10",x"F8",x"4C",x"16",x"82",x"AD",x"FB",x"BC",x"4C",x"24",x"82",x"4C",x"7F",x"8F",x"20",x"34",x"99",x"4C",x"AC",x"8C",x"AE",x"41",x"D6",x"20",x"D0",x"92",x"4C",x"AC",x"8C",x"20",x"98",x"93",x"90",x"03",x"4C",x"16",x"82",x"AD",x"FB",x"BC",x"4C",x"24",x"82",x"20",x"CA",x"93",x"90",x"03",x"4C",x"10",x"82",x"AD",x"FB",x"BC",x"4C",x"24",x"82",x"AE",x"41",x"D6",x"8E",x"F8",x"BC",x"20",x"0D",x"97",x"90",x"0B",x"8D",x"F9",x"BC",x"20",x"84",x"93",x"90",x"03",x"4C",x"16",x"82",x"AD",x"FB",x"BC",x"4C",x"24",x"82",x"20",x"DE",x"93",x"4C",x"AC",x"8C",x"20",x"EB",x"93",x"90",x"03",x"4C",x"10",x"82",x"4C",x"24",x"82",x"20",x"F6",x"93",x"4C",x"AC",x"8C",x"AD",x"FB",x"BC",x"8D",x"40",x"D6",x"4C",x"16",x"82",x"20",x"CE",x"99",x"4C",x"AC",x"8C",x"20",x"4F",x"9A",x"4C",x"AC",x"8C",x"20",x"BC",x"99",x"4C",x"16",x"82",x"20",x"E6",x"8F",x"4C",x"AC",x"8C",x"20",x"A6",x"AB",x"90",x"0B",x"A0",x"00",x"B9",x"00",x"BD",x"91",x"06",x"C8",x"D0",x"F8",x"38",x"4C",x"AC",x"8C",x"AD",x"8B",x"D6",x"29",x"03",x"C9",x"03",x"D0",x"0C",x"09",x"04",x"8D",x"8B",x"D6",x"AD",x"11",x"BD",x"09",x"04",x"38",x"60",x"A9",x"80",x"8D",x"FB",x"BC",x"18",x"60",x"4C",x"35",x"82",x"A9",x"FF",x"8D",x"80",x"BD",x"8D",x"A0",x"BD",x"8D",x"C0",x"BD",x"8D",x"E0",x"BD",x"8D",x"B8",x"BC",x"8D",x"C8",x"BC",x"8D",x"D8",x"BC",x"8D",x"E8",x"BC",x"38",x"60",x"A9",x"00",x"8D",x"FB",x"BC",x"20",x"94",x"90",x"20",x"7D",x"90",x"90",x"3E",x"20",x"BE",x"A0",x"A9",x"02",x"8D",x"FB",x"BC",x"AD",x"FE",x"DF",x"C9",x"55",x"D0",x"2F",x"AD",x"FF",x"DF",x"C9",x"AA",x"D0",x"28",x"A9",x"BE",x"85",x"00",x"A9",x"DF",x"85",x"01",x"20",x"9A",x"90",x"20",x"7D",x"90",x"90",x"18",x"A9",x"CE",x"85",x"00",x"20",x"9A",x"90",x"20",x"7D",x"90",x"90",x"0C",x"A9",x"DE",x"85",x"00",x"20",x"9A",x"90",x"20",x"7D",x"90",x"B0",x"03",x"4C",x"18",x"91",x"A9",x"EE",x"85",x"00",x"20",x"9A",x"90",x"A9",x"00",x"8D",x"FB",x"BC",x"38",x"60",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"82",x"D6",x"8D",x"83",x"D6",x"8D",x"84",x"D6",x"20",x"D3",x"A0",x"B0",x"03",x"4C",x"18",x"91",x"60",x"A9",x"00",x"8D",x"01",x"BC",x"60",x"A9",x"00",x"8D",x"FB",x"BC",x"A0",x"04",x"B1",x"00",x"C9",x"0C",x"F0",x"2C",x"C9",x"0B",x"F0",x"2B",x"C9",x"41",x"F0",x"08",x"A9",x"01",x"8D",x"FB",x"BC",x"4C",x"16",x"91",x"AD",x"FD",x"BC",x"F0",x"03",x"4C",x"18",x"91",x"A0",x"08",x"A2",x"00",x"B1",x"00",x"9D",x"C0",x"BB",x"E8",x"C8",x"C0",x"10",x"D0",x"F5",x"20",x"5E",x"82",x"38",x"60",x"4C",x"D9",x"90",x"4C",x"D9",x"90",x"AD",x"01",x"BC",x"C9",x"06",x"D0",x"03",x"4C",x"18",x"91",x"AD",x"01",x"BC",x"0A",x"0A",x"0A",x"0A",x"0A",x"AA",x"A0",x"08",x"B1",x"00",x"9D",x"00",x"BB",x"E8",x"C8",x"C0",x"10",x"D0",x"F5",x"20",x"1A",x"91",x"90",x"1A",x"AD",x"01",x"BC",x"F0",x"06",x"A0",x"00",x"B1",x"00",x"10",x"08",x"AD",x"01",x"BC",x"8D",x"02",x"BC",x"38",x"60",x"AE",x"01",x"BC",x"38",x"60",x"38",x"60",x"18",x"60",x"A9",x"00",x"8D",x"FB",x"BC",x"AD",x"01",x"BC",x"0A",x"0A",x"0A",x"0A",x"0A",x"8D",x"04",x"BC",x"09",x"00",x"A8",x"A2",x"00",x"B9",x"00",x"BB",x"9D",x"81",x"D6",x"C8",x"E8",x"E0",x"04",x"D0",x"F4",x"20",x"D3",x"A0",x"90",x"D8",x"20",x"BE",x"A0",x"A9",x"02",x"8D",x"FB",x"BC",x"AD",x"FE",x"DF",x"C9",x"55",x"F0",x"03",x"4C",x"18",x"91",x"AD",x"FF",x"DF",x"C9",x"AA",x"F0",x"03",x"4C",x"18",x"91",x"A9",x"03",x"8D",x"FB",x"BC",x"AD",x"11",x"DE",x"D0",x"B2",x"AD",x"04",x"BC",x"09",x"17",x"A8",x"AD",x"10",x"DE",x"99",x"00",x"BB",x"AD",x"04",x"BC",x"09",x"0D",x"A8",x"A2",x"00",x"BD",x"0E",x"DE",x"99",x"00",x"BB",x"C8",x"E8",x"E0",x"02",x"D0",x"F4",x"AD",x"04",x"BC",x"09",x"09",x"A8",x"A2",x"00",x"BD",x"24",x"DE",x"99",x"00",x"BB",x"C8",x"E8",x"E0",x"04",x"D0",x"F4",x"A9",x"04",x"8D",x"FB",x"BC",x"AD",x"2D",x"DE",x"0D",x"2E",x"DE",x"0D",x"2F",x"DE",x"F0",x"03",x"4C",x"18",x"91",x"AC",x"04",x"BC",x"AD",x"2C",x"DE",x"99",x"0F",x"BB",x"AD",x"04",x"BC",x"09",x"0D",x"A8",x"AD",x"04",x"BC",x"09",x"18",x"AA",x"A3",x"02",x"B9",x"00",x"BB",x"9D",x"00",x"BB",x"C8",x"E8",x"3B",x"D0",x"F5",x"6B",x"9D",x"00",x"BB",x"9D",x"01",x"BB",x"A9",x"05",x"8D",x"FB",x"BC",x"AB",x"10",x"DE",x"F0",x"04",x"C2",x"02",x"F0",x"03",x"4C",x"18",x"91",x"AD",x"04",x"BC",x"09",x"18",x"A8",x"A2",x"00",x"18",x"08",x"28",x"B9",x"00",x"BB",x"7D",x"24",x"DE",x"99",x"00",x"BB",x"08",x"C8",x"E8",x"E0",x"04",x"D0",x"EF",x"28",x"3B",x"D0",x"E1",x"AD",x"04",x"BC",x"09",x"18",x"AA",x"AD",x"04",x"BC",x"09",x"12",x"A8",x"38",x"AD",x"20",x"DE",x"FD",x"00",x"BB",x"99",x"00",x"BB",x"AD",x"21",x"DE",x"FD",x"01",x"BB",x"99",x"01",x"BB",x"AD",x"22",x"DE",x"FD",x"02",x"BB",x"99",x"02",x"BB",x"AD",x"23",x"DE",x"FD",x"03",x"BB",x"99",x"03",x"BB",x"AD",x"04",x"BC",x"09",x"16",x"A8",x"AD",x"0D",x"DE",x"99",x"00",x"BB",x"AD",x"0D",x"DE",x"4B",x"29",x"FE",x"F0",x"1E",x"AD",x"04",x"BC",x"09",x"12",x"18",x"69",x"03",x"A8",x"A2",x"03",x"18",x"B9",x"00",x"BB",x"6A",x"99",x"00",x"BB",x"88",x"CA",x"10",x"F5",x"6B",x"4A",x"4B",x"29",x"FE",x"D0",x"E2",x"AD",x"04",x"BC",x"09",x"16",x"A8",x"AD",x"0D",x"DE",x"99",x"00",x"BB",x"AD",x"04",x"BC",x"09",x"16",x"A8",x"A9",x"06",x"8D",x"FB",x"BC",x"B9",x"03",x"BB",x"19",x"02",x"BB",x"D0",x"03",x"4C",x"18",x"91",x"AD",x"04",x"BC",x"09",x"10",x"A8",x"A2",x"03",x"BD",x"2C",x"DE",x"99",x"00",x"BB",x"CA",x"10",x"F7",x"AD",x"04",x"BC",x"09",x"08",x"A8",x"A9",x"0F",x"99",x"00",x"BB",x"EE",x"01",x"BC",x"A9",x"00",x"8D",x"FB",x"BC",x"38",x"60",x"8D",x"FB",x"BC",x"18",x"60",x"EC",x"01",x"BC",x"90",x"07",x"A9",x"80",x"8D",x"FB",x"BC",x"18",x"60",x"8E",x"03",x"BC",x"8A",x"0A",x"0A",x"0A",x"0A",x"0A",x"8D",x"04",x"BC",x"38",x"60",x"20",x"B6",x"92",x"B0",x"02",x"18",x"60",x"AE",x"04",x"BC",x"BD",x"10",x"BB",x"8D",x"05",x"BC",x"BD",x"11",x"BB",x"8D",x"06",x"BC",x"A9",x"00",x"8D",x"07",x"BC",x"8D",x"08",x"BC",x"4C",x"AA",x"92",x"A2",x"03",x"BD",x"B3",x"BC",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"A9",x"FF",x"AA",x"A8",x"4B",x"A9",x"FE",x"20",x"0B",x"9C",x"AE",x"04",x"BC",x"BD",x"16",x"BB",x"A8",x"29",x"FE",x"F0",x"14",x"18",x"2E",x"81",x"D6",x"2E",x"82",x"D6",x"2E",x"83",x"D6",x"2E",x"84",x"D6",x"98",x"4A",x"A8",x"29",x"FE",x"D0",x"EC",x"A9",x"18",x"20",x"2A",x"9C",x"A9",x"00",x"20",x"2A",x"9C",x"38",x"60",x"A2",x"00",x"8A",x"0A",x"0A",x"0A",x"0A",x"A8",x"B9",x"B8",x"BC",x"C9",x"FF",x"F0",x"0A",x"E8",x"E0",x"04",x"D0",x"EE",x"A9",x"84",x"4C",x"B1",x"92",x"8E",x"F8",x"BC",x"8C",x"F9",x"BC",x"18",x"A9",x"B8",x"6D",x"F9",x"BC",x"A8",x"A9",x"BC",x"69",x"00",x"48",x"5A",x"A0",x"0F",x"A9",x"00",x"82",x"01",x"88",x"D0",x"FB",x"68",x"68",x"38",x"60",x"A9",x"FF",x"8D",x"B8",x"BC",x"8D",x"C8",x"BC",x"8D",x"D8",x"BC",x"8D",x"E8",x"BC",x"A2",x"00",x"A9",x"00",x"9D",x"00",x"BB",x"E8",x"D0",x"FA",x"38",x"60",x"AE",x"F9",x"BC",x"BD",x"B9",x"BC",x"C9",x"01",x"D0",x"00",x"AE",x"F9",x"BC",x"A9",x"FF",x"9D",x"B8",x"BC",x"38",x"60",x"AD",x"65",x"BC",x"29",x"10",x"D0",x"05",x"A9",x"87",x"4C",x"B1",x"92",x"20",x"99",x"96",x"90",x"47",x"20",x"84",x"93",x"A2",x"03",x"BD",x"5D",x"BC",x"9D",x"05",x"BC",x"CA",x"10",x"F7",x"A2",x"03",x"A9",x"00",x"1D",x"05",x"BC",x"CA",x"10",x"FA",x"C9",x"00",x"D0",x"03",x"4C",x"D7",x"92",x"38",x"60",x"AD",x"65",x"BC",x"29",x"10",x"F0",x"05",x"A9",x"86",x"4C",x"B1",x"92",x"20",x"99",x"96",x"90",x"15",x"4C",x"E6",x"96",x"20",x"EB",x"93",x"B0",x"03",x"4C",x"F0",x"93",x"20",x"84",x"93",x"38",x"60",x"20",x"0A",x"94",x"B0",x"03",x"4C",x"B4",x"92",x"4C",x"F6",x"93",x"20",x"45",x"94",x"B0",x"08",x"20",x"84",x"93",x"A9",x"88",x"4C",x"B1",x"92",x"20",x"52",x"96",x"90",x"EE",x"38",x"60",x"A9",x"80",x"0C",x"89",x"D6",x"20",x"31",x"93",x"B0",x"03",x"4C",x"B4",x"92",x"8A",x"0A",x"0A",x"0A",x"0A",x"A8",x"AD",x"03",x"BC",x"99",x"B8",x"BC",x"A2",x"00",x"BD",x"05",x"BC",x"99",x"BA",x"BC",x"99",x"BE",x"BC",x"C8",x"E8",x"E0",x"04",x"D0",x"F1",x"AE",x"F9",x"BC",x"A9",x"80",x"9D",x"B9",x"BC",x"20",x"E6",x"96",x"B0",x"03",x"4C",x"B4",x"92",x"60",x"A9",x"00",x"8D",x"4F",x"BC",x"AE",x"F9",x"BC",x"BD",x"B9",x"BC",x"C9",x"81",x"D0",x"05",x"A9",x"FF",x"4C",x"B1",x"92",x"20",x"34",x"97",x"AE",x"F9",x"BC",x"BD",x"B9",x"BC",x"C9",x"80",x"F0",x"0E",x"C9",x"81",x"D0",x"05",x"A9",x"FF",x"4C",x"B1",x"92",x"A9",x"87",x"4C",x"B1",x"92",x"A2",x"56",x"A9",x"00",x"9D",x"0F",x"BC",x"CA",x"10",x"FA",x"20",x"34",x"97",x"B0",x"03",x"4C",x"B4",x"92",x"20",x"BE",x"A0",x"AD",x"F9",x"BC",x"09",x"0B",x"AA",x"BD",x"B8",x"BC",x"85",x"00",x"BD",x"B9",x"BC",x"18",x"69",x"DE",x"85",x"01",x"A0",x"00",x"B1",x"00",x"C9",x"E5",x"D0",x"03",x"4C",x"42",x"96",x"C9",x"00",x"D0",x"03",x"4C",x"42",x"96",x"A0",x"0B",x"B1",x"00",x"A8",x"29",x"0F",x"C9",x"0F",x"D0",x"03",x"4C",x"D1",x"94",x"98",x"29",x"08",x"C9",x"08",x"D0",x"03",x"4C",x"6E",x"95",x"98",x"29",x"06",x"F0",x"03",x"4C",x"6E",x"95",x"4C",x"79",x"95",x"4C",x"6E",x"95",x"A0",x"0C",x"B1",x"00",x"F0",x"03",x"4C",x"79",x"95",x"A0",x"00",x"B1",x"00",x"48",x"29",x"40",x"8D",x"FA",x"BC",x"68",x"29",x"3F",x"3A",x"C9",x"05",x"B0",x"72",x"AA",x"BD",x"4D",x"96",x"AA",x"A0",x"01",x"A3",x"05",x"B1",x"00",x"F0",x"58",x"20",x"E7",x"9F",x"9D",x"0F",x"BC",x"AD",x"FA",x"BC",x"F0",x"03",x"8E",x"4F",x"BC",x"E8",x"E0",x"40",x"F0",x"45",x"C8",x"C8",x"3B",x"D0",x"E4",x"A0",x"0E",x"A3",x"06",x"B1",x"00",x"F0",x"38",x"20",x"E7",x"9F",x"9D",x"0F",x"BC",x"AD",x"FA",x"BC",x"F0",x"03",x"8E",x"4F",x"BC",x"E8",x"E0",x"40",x"F0",x"25",x"C8",x"C8",x"3B",x"D0",x"E4",x"A0",x"1C",x"A3",x"02",x"B1",x"00",x"F0",x"18",x"20",x"E7",x"9F",x"9D",x"0F",x"BC",x"AD",x"FA",x"BC",x"F0",x"03",x"8E",x"4F",x"BC",x"E8",x"E0",x"40",x"F0",x"05",x"C8",x"C8",x"3B",x"D0",x"E4",x"AD",x"FA",x"BC",x"F0",x"08",x"EC",x"4F",x"BC",x"90",x"03",x"8E",x"4F",x"BC",x"20",x"70",x"96",x"90",x"03",x"4C",x"89",x"94",x"A9",x"FF",x"4C",x"B1",x"92",x"20",x"70",x"96",x"90",x"03",x"4C",x"45",x"94",x"4C",x"B4",x"92",x"A0",x"00",x"A2",x"00",x"B1",x"00",x"9D",x"50",x"BC",x"E8",x"C8",x"E0",x"0B",x"D0",x"F5",x"AD",x"4F",x"BC",x"D0",x"5B",x"A0",x"00",x"A2",x"00",x"B1",x"00",x"9D",x"0F",x"BC",x"8E",x"4F",x"BC",x"E8",x"C8",x"C9",x"20",x"F0",x"05",x"E0",x"08",x"D0",x"EE",x"E8",x"CA",x"A9",x"2E",x"9D",x"0F",x"BC",x"8E",x"4F",x"BC",x"E8",x"A0",x"08",x"A3",x"00",x"B1",x"00",x"9D",x"0F",x"BC",x"8E",x"4F",x"BC",x"E8",x"C8",x"1B",x"C2",x"03",x"F0",x"08",x"C9",x"20",x"F0",x"04",x"E0",x"0C",x"D0",x"E9",x"E0",x"00",x"F0",x"13",x"A9",x"20",x"DD",x"0E",x"BC",x"D0",x"04",x"CA",x"4C",x"C9",x"95",x"BD",x"0E",x"BC",x"C9",x"2E",x"D0",x"01",x"CA",x"A9",x"00",x"9D",x"0F",x"BC",x"8E",x"4F",x"BC",x"A0",x"1A",x"B1",x"00",x"8D",x"5D",x"BC",x"C8",x"B1",x"00",x"8D",x"5E",x"BC",x"A0",x"14",x"B1",x"00",x"8D",x"5F",x"BC",x"C8",x"B1",x"00",x"8D",x"60",x"BC",x"A0",x"1C",x"A2",x"00",x"B1",x"00",x"9D",x"61",x"BC",x"C8",x"E8",x"E0",x"04",x"D0",x"F5",x"A0",x"0B",x"B1",x"00",x"8D",x"65",x"BC",x"20",x"70",x"96",x"B0",x"10",x"AE",x"F9",x"BC",x"A9",x"81",x"9D",x"B9",x"BC",x"AE",x"F9",x"BC",x"BD",x"B9",x"BC",x"38",x"60",x"AD",x"4F",x"BC",x"C9",x"00",x"F0",x"09",x"AD",x"50",x"BC",x"F0",x"04",x"C9",x"20",x"D0",x"03",x"4C",x"45",x"94",x"38",x"60",x"20",x"70",x"96",x"90",x"03",x"4C",x"45",x"94",x"4C",x"B4",x"92",x"00",x"0D",x"1A",x"27",x"34",x"AD",x"4F",x"BC",x"CD",x"66",x"BC",x"D0",x"14",x"AE",x"4F",x"BC",x"CA",x"BD",x"67",x"BC",x"20",x"E7",x"9F",x"DD",x"0F",x"BC",x"D0",x"05",x"CA",x"10",x"F2",x"38",x"60",x"18",x"60",x"AC",x"F9",x"BC",x"18",x"B9",x"C3",x"BC",x"69",x"20",x"99",x"C3",x"BC",x"D0",x"0B",x"B9",x"C4",x"BC",x"1A",x"C9",x"01",x"D0",x"05",x"99",x"C4",x"BC",x"38",x"60",x"A9",x"00",x"99",x"C4",x"BC",x"20",x"51",x"97",x"90",x"03",x"20",x"34",x"97",x"60",x"20",x"31",x"93",x"20",x"0D",x"97",x"B0",x"03",x"4C",x"B4",x"92",x"AD",x"03",x"BC",x"9D",x"B8",x"BC",x"A0",x"00",x"B9",x"5D",x"BC",x"9D",x"BA",x"BC",x"9D",x"BE",x"BC",x"E8",x"C8",x"C0",x"04",x"D0",x"F1",x"20",x"0D",x"97",x"B0",x"03",x"4C",x"B4",x"92",x"AD",x"03",x"BC",x"9D",x"B8",x"BC",x"A9",x"00",x"9D",x"B9",x"BC",x"A9",x"00",x"9D",x"C2",x"BC",x"9D",x"C3",x"BC",x"9D",x"C4",x"BC",x"A2",x"03",x"BD",x"61",x"BC",x"9D",x"AB",x"BC",x"CA",x"10",x"F7",x"38",x"60",x"20",x"0D",x"97",x"B0",x"03",x"4C",x"B4",x"92",x"A0",x"03",x"BD",x"BA",x"BC",x"9D",x"BE",x"BC",x"E8",x"88",x"10",x"F6",x"20",x"0D",x"97",x"A9",x"00",x"A0",x"06",x"9D",x"C2",x"BC",x"E8",x"88",x"D0",x"F9",x"20",x"0D",x"97",x"38",x"60",x"AD",x"F8",x"BC",x"C9",x"04",x"B0",x"07",x"0A",x"0A",x"0A",x"0A",x"AA",x"38",x"60",x"A9",x"89",x"4C",x"B1",x"92",x"20",x"0D",x"97",x"90",x"1D",x"A0",x"00",x"BD",x"BE",x"BC",x"99",x"B3",x"BC",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"60",x"20",x"0D",x"97",x"20",x"20",x"97",x"20",x"F1",x"92",x"20",x"0D",x"97",x"B0",x"03",x"4C",x"B4",x"92",x"09",x"0A",x"A8",x"B9",x"B8",x"BC",x"20",x"04",x"9C",x"4C",x"D3",x"A0",x"AE",x"F9",x"BC",x"BD",x"C5",x"BC",x"18",x"69",x"02",x"9D",x"C5",x"BC",x"90",x"08",x"FE",x"C6",x"BC",x"D0",x"03",x"FE",x"C7",x"BC",x"FE",x"C2",x"BC",x"BD",x"C2",x"BC",x"AC",x"04",x"BC",x"D9",x"16",x"BB",x"F0",x"02",x"38",x"60",x"AC",x"F9",x"BC",x"A9",x"00",x"99",x"C2",x"BC",x"20",x"20",x"97",x"A2",x"03",x"BD",x"B3",x"BC",x"9D",x"AF",x"BC",x"CA",x"10",x"F7",x"AD",x"B3",x"BC",x"8D",x"04",x"BF",x"20",x"54",x"98",x"20",x"39",x"98",x"A2",x"03",x"08",x"BD",x"B3",x"BC",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"28",x"BD",x"B3",x"BC",x"69",x"00",x"9D",x"B3",x"BC",x"08",x"E8",x"E0",x"04",x"D0",x"F1",x"28",x"20",x"D3",x"A0",x"B0",x"03",x"4C",x"B4",x"92",x"20",x"BE",x"A0",x"AD",x"04",x"BF",x"0A",x"0A",x"AA",x"AD",x"F9",x"BC",x"09",x"06",x"A8",x"8C",x"05",x"BF",x"AC",x"05",x"BF",x"A3",x"00",x"AD",x"04",x"BF",x"29",x"40",x"D0",x"0F",x"BD",x"00",x"DE",x"99",x"B8",x"BC",x"E8",x"C8",x"1B",x"C2",x"04",x"D0",x"F3",x"80",x"0D",x"BD",x"00",x"DF",x"99",x"B8",x"BC",x"E8",x"C8",x"1B",x"C2",x"04",x"D0",x"F3",x"AC",x"05",x"BF",x"B9",x"BB",x"BC",x"29",x"0F",x"99",x"BB",x"BC",x"B9",x"BB",x"BC",x"19",x"BA",x"BC",x"19",x"B9",x"BC",x"19",x"B8",x"BC",x"C9",x"00",x"F0",x"1F",x"B9",x"BB",x"BC",x"C9",x"0F",x"D0",x"13",x"B9",x"BA",x"BC",x"39",x"B9",x"BC",x"C9",x"FF",x"D0",x"09",x"B9",x"B8",x"BC",x"29",x"F0",x"C9",x"F0",x"F0",x"05",x"20",x"45",x"98",x"38",x"60",x"20",x"45",x"98",x"A9",x"85",x"4C",x"B1",x"92",x"A2",x"03",x"BD",x"81",x"D6",x"9D",x"55",x"BD",x"CA",x"10",x"F7",x"60",x"A2",x"03",x"BD",x"55",x"BD",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"20",x"D3",x"A0",x"60",x"A0",x"07",x"18",x"6E",x"B6",x"BC",x"6E",x"B5",x"BC",x"6E",x"B4",x"BC",x"6E",x"B3",x"BC",x"88",x"D0",x"F0",x"AC",x"04",x"BC",x"A2",x"00",x"18",x"08",x"28",x"BD",x"B3",x"BC",x"79",x"00",x"BB",x"9D",x"B3",x"BC",x"08",x"C8",x"E8",x"E0",x"04",x"D0",x"EF",x"28",x"AC",x"04",x"BC",x"A2",x"00",x"18",x"08",x"28",x"BD",x"B3",x"BC",x"79",x"0D",x"BB",x"9D",x"B3",x"BC",x"08",x"C8",x"E8",x"E0",x"02",x"D0",x"EF",x"28",x"60",x"A2",x"00",x"8E",x"A9",x"BC",x"8E",x"AA",x"BC",x"20",x"EB",x"93",x"90",x"0E",x"20",x"84",x"93",x"20",x"CA",x"93",x"90",x"06",x"20",x"BE",x"A0",x"4C",x"B7",x"98",x"4C",x"B4",x"92",x"20",x"34",x"97",x"90",x"3D",x"20",x"FF",x"98",x"A2",x"00",x"A3",x"00",x"BD",x"00",x"DE",x"EA",x"92",x"18",x"1B",x"E8",x"88",x"D0",x"F5",x"E3",x"19",x"20",x"FF",x"98",x"BD",x"00",x"DF",x"EA",x"92",x"18",x"1B",x"E8",x"88",x"D0",x"F5",x"20",x"51",x"97",x"90",x"16",x"E3",x"19",x"EE",x"A9",x"BC",x"D0",x"CD",x"EE",x"AA",x"BC",x"D0",x"C8",x"20",x"84",x"93",x"A9",x"83",x"4C",x"B1",x"92",x"68",x"68",x"20",x"84",x"93",x"4C",x"AA",x"92",x"A0",x"00",x"AD",x"AC",x"BC",x"0D",x"AD",x"BC",x"0D",x"AE",x"BC",x"D0",x"0E",x"AD",x"AB",x"BC",x"F0",x"E6",x"AC",x"AB",x"BC",x"A9",x"00",x"8D",x"AB",x"BC",x"60",x"AD",x"AC",x"BC",x"38",x"E9",x"01",x"8D",x"AC",x"BC",x"AD",x"AD",x"BC",x"E9",x"00",x"8D",x"AD",x"BC",x"AD",x"AE",x"BC",x"E9",x"00",x"8D",x"AE",x"BC",x"60",x"AD",x"AB",x"BC",x"0D",x"AC",x"BC",x"0D",x"AD",x"BC",x"0D",x"AE",x"BC",x"D0",x"0A",x"A9",x"00",x"8D",x"41",x"D6",x"8D",x"42",x"D6",x"18",x"60",x"A2",x"00",x"A0",x"02",x"AD",x"AD",x"BC",x"0D",x"AE",x"BC",x"D0",x"17",x"AD",x"AC",x"BC",x"C9",x"02",x"B0",x"10",x"AE",x"AB",x"BC",x"AC",x"AC",x"BC",x"A9",x"00",x"8D",x"AB",x"BC",x"A9",x"02",x"8D",x"AC",x"BC",x"AD",x"AC",x"BC",x"38",x"E9",x"02",x"8D",x"AC",x"BC",x"AD",x"AD",x"BC",x"E9",x"00",x"8D",x"AD",x"BC",x"AD",x"AE",x"BC",x"E9",x"00",x"8D",x"AE",x"BC",x"8E",x"41",x"D6",x"8C",x"42",x"D6",x"20",x"BE",x"A0",x"20",x"34",x"97",x"B0",x"01",x"60",x"20",x"51",x"97",x"38",x"60",x"86",x"00",x"84",x"01",x"A0",x"00",x"B1",x"00",x"99",x"67",x"BC",x"F0",x"0E",x"C8",x"C0",x"40",x"D0",x"F4",x"A9",x"00",x"8D",x"66",x"BC",x"A9",x"81",x"18",x"60",x"8C",x"66",x"BC",x"38",x"60",x"A9",x"00",x"8D",x"8B",x"D6",x"8D",x"8A",x"D6",x"A9",x"01",x"1C",x"11",x"BD",x"1C",x"12",x"BD",x"38",x"60",x"20",x"DE",x"93",x"B0",x"04",x"A9",x"88",x"18",x"60",x"20",x"84",x"93",x"20",x"D0",x"9A",x"B0",x"01",x"60",x"A2",x"03",x"BD",x"81",x"D6",x"9D",x"8C",x"D6",x"CA",x"10",x"F7",x"AD",x"A1",x"D6",x"29",x"FE",x"8D",x"A1",x"D6",x"AD",x"8B",x"D6",x"29",x"B8",x"09",x"07",x"8D",x"8B",x"D6",x"A9",x"40",x"1C",x"8A",x"D6",x"AD",x"27",x"BF",x"C9",x"40",x"D0",x"08",x"A9",x"40",x"0C",x"8A",x"D6",x"4C",x"29",x"9A",x"C9",x"47",x"D0",x"0B",x"A9",x"40",x"0C",x"8A",x"D6",x"0C",x"8B",x"D6",x"4C",x"29",x"9A",x"C9",x"41",x"D0",x"05",x"A9",x"40",x"0C",x"8B",x"D6",x"A9",x"01",x"8D",x"11",x"BD",x"AE",x"66",x"BC",x"E0",x"20",x"B0",x"13",x"8E",x"13",x"BD",x"A2",x"00",x"BD",x"67",x"BC",x"9D",x"15",x"BD",x"E8",x"EC",x"13",x"BD",x"D0",x"F4",x"38",x"60",x"A9",x"00",x"8D",x"13",x"BD",x"38",x"60",x"20",x"DE",x"93",x"B0",x"04",x"A9",x"88",x"18",x"60",x"20",x"84",x"93",x"20",x"D0",x"9A",x"B0",x"01",x"60",x"A2",x"03",x"BD",x"81",x"D6",x"9D",x"90",x"D6",x"CA",x"10",x"F7",x"AD",x"A1",x"D6",x"29",x"FB",x"8D",x"A1",x"D6",x"AD",x"8B",x"D6",x"29",x"47",x"09",x"38",x"8D",x"8B",x"D6",x"A9",x"80",x"1C",x"8A",x"D6",x"AD",x"27",x"BF",x"C9",x"40",x"D0",x"08",x"A9",x"80",x"0C",x"8A",x"D6",x"4C",x"AA",x"9A",x"C9",x"47",x"D0",x"0B",x"A9",x"80",x"0C",x"8A",x"D6",x"0C",x"8B",x"D6",x"4C",x"AA",x"9A",x"C9",x"41",x"D0",x"05",x"A9",x"80",x"0C",x"8B",x"D6",x"A9",x"01",x"8D",x"12",x"BD",x"AE",x"66",x"BC",x"E0",x"20",x"B0",x"13",x"8E",x"14",x"BD",x"A2",x"00",x"BD",x"67",x"BC",x"9D",x"35",x"BD",x"E8",x"EC",x"14",x"BD",x"D0",x"F4",x"38",x"60",x"A9",x"00",x"8D",x"14",x"BD",x"38",x"60",x"20",x"99",x"96",x"90",x"05",x"20",x"CA",x"93",x"B0",x"03",x"4C",x"02",x"9C",x"A9",x"00",x"8D",x"32",x"BF",x"8D",x"33",x"BF",x"A9",x"40",x"8D",x"2C",x"BF",x"A9",x"06",x"8D",x"2D",x"BF",x"A9",x"58",x"8D",x"2E",x"BF",x"A9",x"01",x"8D",x"2F",x"BF",x"A9",x"B0",x"8D",x"30",x"BF",x"A9",x"02",x"8D",x"31",x"BF",x"AE",x"04",x"BC",x"BD",x"16",x"BB",x"4B",x"6B",x"29",x"01",x"D0",x"18",x"6B",x"4A",x"4B",x"4E",x"2D",x"BF",x"6E",x"2C",x"BF",x"4E",x"2F",x"BF",x"6E",x"2E",x"BF",x"4E",x"31",x"BF",x"6E",x"30",x"BF",x"4C",x"0A",x"9B",x"AE",x"F9",x"BC",x"A0",x"00",x"BD",x"BE",x"BC",x"99",x"28",x"BF",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"AE",x"F9",x"BC",x"A0",x"00",x"BD",x"BE",x"BC",x"D9",x"28",x"BF",x"F0",x"03",x"4C",x"F8",x"9B",x"E8",x"C8",x"C0",x"04",x"D0",x"EF",x"EE",x"32",x"BF",x"D0",x"03",x"EE",x"33",x"BF",x"18",x"AD",x"28",x"BF",x"69",x"01",x"8D",x"28",x"BF",x"AD",x"29",x"BF",x"69",x"00",x"8D",x"29",x"BF",x"AD",x"2A",x"BF",x"69",x"00",x"8D",x"2A",x"BF",x"AD",x"2B",x"BF",x"69",x"00",x"8D",x"2B",x"BF",x"20",x"77",x"97",x"B0",x"BC",x"A9",x"00",x"8D",x"FB",x"BC",x"20",x"84",x"93",x"AD",x"34",x"BF",x"0D",x"35",x"BF",x"D0",x"65",x"AD",x"33",x"BF",x"CD",x"2F",x"BF",x"D0",x"0F",x"AD",x"32",x"BF",x"CD",x"2E",x"BF",x"D0",x"04",x"A9",x"40",x"80",x"38",x"AD",x"33",x"BF",x"CD",x"31",x"BF",x"D0",x"0F",x"AD",x"32",x"BF",x"CD",x"30",x"BF",x"D0",x"04",x"A9",x"47",x"80",x"24",x"AD",x"33",x"BF",x"C9",x"05",x"D0",x"0E",x"AD",x"32",x"BF",x"C9",x"50",x"D0",x"04",x"A9",x"41",x"80",x"12",x"AD",x"2D",x"BF",x"CD",x"33",x"BF",x"D0",x"23",x"AD",x"2C",x"BF",x"CD",x"32",x"BF",x"D0",x"1B",x"A9",x"51",x"8D",x"27",x"BF",x"AE",x"F9",x"BC",x"A0",x"00",x"BD",x"BA",x"BC",x"99",x"B3",x"BC",x"E8",x"C8",x"C0",x"04",x"D0",x"F4",x"20",x"F1",x"92",x"38",x"60",x"A9",x"8A",x"8D",x"FB",x"BC",x"18",x"60",x"20",x"84",x"93",x"A9",x"8B",x"8D",x"FB",x"BC",x"18",x"60",x"18",x"60",x"48",x"A9",x"00",x"AA",x"A8",x"4B",x"68",x"18",x"6D",x"81",x"D6",x"8D",x"81",x"D6",x"8A",x"6D",x"82",x"D6",x"8D",x"82",x"D6",x"98",x"6D",x"83",x"D6",x"8D",x"83",x"D6",x"6B",x"6D",x"84",x"D6",x"8D",x"84",x"D6",x"A3",x"00",x"60",x"0D",x"04",x"BC",x"A8",x"A2",x"00",x"18",x"08",x"28",x"BD",x"81",x"D6",x"79",x"00",x"BB",x"9D",x"81",x"D6",x"08",x"C8",x"E8",x"E0",x"04",x"D0",x"EF",x"28",x"60",x"C9",x"20",x"90",x"05",x"C9",x"7F",x"B0",x"01",x"60",x"A9",x"3F",x"60",x"20",x"BE",x"A0",x"A9",x"02",x"8D",x"09",x"BC",x"8D",x"18",x"BF",x"A9",x"00",x"8D",x"0A",x"BC",x"8D",x"0B",x"BC",x"8D",x"0C",x"BC",x"8D",x"19",x"BF",x"8D",x"1A",x"BF",x"8D",x"1B",x"BF",x"A2",x"03",x"BD",x"61",x"BC",x"9D",x"5D",x"BC",x"CA",x"10",x"F7",x"A2",x"03",x"BD",x"18",x"BF",x"9D",x"B3",x"BC",x"CA",x"10",x"F7",x"20",x"54",x"98",x"A2",x"03",x"BD",x"B3",x"BC",x"9D",x"81",x"D6",x"CA",x"10",x"F7",x"A9",x"20",x"8D",x"FB",x"BC",x"20",x"D3",x"A0",x"B0",x"01",x"60",x"AE",x"03",x"BC",x"20",x"B6",x"92",x"AE",x"04",x"BC",x"A0",x"00",x"BD",x"12",x"BB",x"D9",x"18",x"BF",x"D0",x"0D",x"E8",x"C8",x"C0",x"04",x"D0",x"F2",x"A9",x"8C",x"8D",x"FB",x"BC",x"18",x"60",x"AD",x"18",x"BF",x"0A",x"0A",x"A8",x"AD",x"18",x"BF",x"29",x"40",x"F0",x"0E",x"B9",x"00",x"DF",x"19",x"01",x"DF",x"19",x"02",x"DF",x"19",x"03",x"DF",x"80",x"0C",x"B9",x"00",x"DE",x"19",x"01",x"DE",x"19",x"02",x"DE",x"19",x"03",x"DE",x"AA",x"AD",x"18",x"BF",x"18",x"69",x"01",x"8D",x"18",x"BF",x"AD",x"19",x"BF",x"69",x"00",x"AD",x"19",x"BF",x"AD",x"1A",x"BF",x"69",x"00",x"AD",x"1A",x"BF",x"AD",x"1B",x"BF",x"69",x"00",x"AD",x"1B",x"BF",x"E0",x"00",x"F0",x"0E",x"A2",x"03",x"BD",x"18",x"BF",x"9D",x"09",x"BC",x"CA",x"10",x"F7",x"4C",x"70",x"9C",x"AD",x"5D",x"BC",x"38",x"E9",x"01",x"8D",x"5D",x"BC",x"AD",x"5E",x"BC",x"E9",x"00",x"8D",x"5E",x"BC",x"AD",x"5F",x"BC",x"E9",x"00",x"8D",x"5F",x"BC",x"AD",x"60",x"BC",x"E9",x"00",x"8D",x"60",x"BC",x"0D",x"5F",x"BC",x"0D",x"5E",x"BC",x"0D",x"5D",x"BC",x"F0",x"0D",x"AD",x"18",x"BF",x"29",x"7F",x"D0",x"03",x"4C",x"7B",x"9C",x"4C",x"9F",x"9C",x"38",x"60",x"20",x"45",x"A3",x"A2",x"85",x"A0",x"9D",x"20",x"2B",x"A9",x"A0",x"00",x"AB",x"49",x"D6",x"20",x"A4",x"A9",x"AB",x"48",x"D6",x"20",x"A4",x"A9",x"AB",x"4F",x"D6",x"20",x"A4",x"A9",x"AB",x"4A",x"D6",x"20",x"A4",x"A9",x"AB",x"49",x"D6",x"20",x"A4",x"A9",x"EE",x"20",x"D0",x"4C",x"7F",x"9D",x"50",x"41",x"47",x"45",x"20",x"46",x"41",x"55",x"4C",x"54",x"3A",x"20",x"50",x"43",x"3D",x"24",x"24",x"24",x"24",x"2C",x"20",x"4D",x"41",x"50",x"3D",x"24",x"24",x"2E",x"24",x"24",x"24",x"24",x"2E",x"30",x"30",x"20",x"20",x"20",x"20",x"20",x"78",x"D8",x"29",x"FE",x"AA",x"7C",x"B5",x"9D",x"3D",x"9E",x"35",x"9E",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"35",x"82",x"A9",x"04",x"1C",x"7D",x"D6",x"4C",x"16",x"82",x"A9",x"04",x"0C",x"7D",x"D6",x"4C",x"16",x"82",x"A9",x"00",x"60",x"A9",x"00",x"8D",x"40",x"D6",x"8D",x"41",x"D6",x"8D",x"42",x"D6",x"8D",x"43",x"D6",x"8D",x"44",x"D6",x"A9",x"FF",x"8D",x"45",x"D6",x"A9",x"01",x"8D",x"46",x"D6",x"A9",x"F7",x"8D",x"47",x"D6",x"A9",x"00",x"8D",x"4A",x"D6",x"8D",x"4B",x"D6",x"8D",x"4C",x"D6",x"8D",x"4D",x"D6",x"8D",x"4E",x"D6",x"8D",x"4F",x"D6",x"A9",x"3F",x"8D",x"50",x"D6",x"8D",x"51",x"D6",x"A9",x"00",x"8D",x"52",x"D6",x"A9",x"82",x"8D",x"80",x"D6",x"A9",x"01",x"1C",x"30",x"D0",x"A9",x"D7",x"1C",x"54",x"D0",x"A9",x"00",x"8D",x"30",x"D0",x"8D",x"31",x"D0",x"AD",x"00",x"DD",x"09",x"03",x"8D",x"00",x"DD",x"A9",x"C0",x"8D",x"5D",x"D0",x"A9",x"1B",x"8D",x"11",x"D0",x"A9",x"C8",x"8D",x"16",x"D0",x"A9",x"14",x"8D",x"18",x"D0",x"60",x"A2",x"FC",x"A0",x"FF",x"A3",x"02",x"A9",x"00",x"20",x"A4",x"AA",x"AD",x"00",x"BC",x"8D",x"48",x"D6",x"A2",x"FC",x"E8",x"A0",x"FF",x"A3",x"02",x"A9",x"00",x"20",x"A4",x"AA",x"AD",x"00",x"BC",x"8D",x"49",x"D6",x"60",x"A9",x"C1",x"8D",x"18",x"03",x"A9",x"FE",x"8D",x"19",x"03",x"60",x"A9",x"00",x"A2",x"5D",x"9D",x"00",x"D6",x"E8",x"E0",x"70",x"D0",x"F8",x"60",x"A2",x"00",x"8A",x"9D",x"00",x"BD",x"E8",x"D0",x"FA",x"20",x"EC",x"9E",x"4C",x"05",x"90",x"20",x"F9",x"9E",x"20",x"45",x"9E",x"8D",x"00",x"BD",x"60",x"20",x"08",x"9F",x"20",x"48",x"9E",x"60",x"A9",x"FF",x"8D",x"00",x"BD",x"60",x"AD",x"00",x"BD",x"C9",x"FF",x"D0",x"03",x"8D",x"7F",x"D6",x"A9",x"01",x"1C",x"30",x"D0",x"A9",x"00",x"8D",x"11",x"D7",x"AA",x"A8",x"20",x"90",x"86",x"20",x"19",x"9F",x"20",x"9F",x"A6",x"20",x"B9",x"A6",x"A2",x"43",x"A0",x"B3",x"20",x"9C",x"99",x"AE",x"02",x"BC",x"20",x"D0",x"92",x"A9",x"00",x"85",x"1A",x"85",x"1B",x"A9",x"07",x"85",x"19",x"A9",x"FF",x"85",x"18",x"20",x"99",x"98",x"EE",x"20",x"D0",x"90",x"F8",x"CE",x"20",x"D0",x"20",x"48",x"9E",x"20",x"E1",x"9E",x"A9",x"0D",x"8D",x"48",x"D6",x"A9",x"08",x"8D",x"49",x"D6",x"A9",x"FF",x"8D",x"26",x"03",x"A9",x"03",x"8D",x"27",x"03",x"A9",x"60",x"8D",x"FF",x"03",x"A9",x"FC",x"8D",x"14",x"03",x"8D",x"16",x"03",x"8D",x"18",x"03",x"A9",x"03",x"8D",x"15",x"03",x"8D",x"17",x"03",x"8D",x"19",x"03",x"A9",x"4C",x"8D",x"FC",x"03",x"A9",x"81",x"8D",x"FD",x"03",x"A9",x"EA",x"8D",x"FE",x"03",x"A9",x"7F",x"8D",x"0D",x"DC",x"8D",x"0D",x"DD",x"A9",x"00",x"8D",x"1A",x"D0",x"8D",x"7F",x"D6",x"AD",x"40",x"D6",x"8D",x"72",x"D6",x"8D",x"7F",x"D6",x"AD",x"72",x"D6",x"49",x"40",x"8D",x"72",x"D6",x"8D",x"7F",x"D6",x"A9",x"32",x"8D",x"7D",x"D6",x"A9",x"C0",x"8D",x"72",x"D6",x"4C",x"00",x"82",x"EE",x"21",x"D0",x"A9",x"00",x"8D",x"72",x"D6",x"4C",x"00",x"82",x"C9",x"61",x"90",x"06",x"C9",x"7B",x"B0",x"02",x"29",x"5F",x"60",x"20",x"6A",x"A0",x"B0",x"01",x"60",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"82",x"D6",x"8D",x"83",x"D6",x"8D",x"84",x"D6",x"A9",x"40",x"8D",x"80",x"D6",x"A9",x"02",x"8D",x"81",x"D6",x"8D",x"80",x"D6",x"20",x"A2",x"A0",x"B0",x"17",x"D0",x"F9",x"A9",x"00",x"8D",x"81",x"D6",x"20",x"6A",x"A0",x"A2",x"4D",x"A0",x"AF",x"20",x"2B",x"A9",x"EE",x"20",x"D0",x"4C",x"29",x"A0",x"A2",x"70",x"A0",x"AF",x"20",x"2B",x"A9",x"A9",x"41",x"8D",x"80",x"D6",x"4C",x"D3",x"A0",x"A9",x"57",x"8D",x"80",x"D6",x"60",x"20",x"3E",x"A0",x"4C",x"4F",x"A0",x"A9",x"4D",x"8D",x"80",x"D6",x"A9",x"03",x"8D",x"80",x"D6",x"60",x"20",x"94",x"A0",x"20",x"A2",x"A0",x"90",x"FB",x"60",x"20",x"55",x"A0",x"B0",x"06",x"20",x"6A",x"A0",x"4C",x"5E",x"A0",x"60",x"A9",x"00",x"8D",x"80",x"D6",x"A9",x"01",x"8D",x"80",x"D6",x"20",x"55",x"A0",x"B0",x"03",x"D0",x"F9",x"60",x"20",x"BE",x"A0",x"38",x"60",x"20",x"94",x"A0",x"EE",x"1C",x"BF",x"D0",x"FB",x"EE",x"1D",x"BF",x"D0",x"F6",x"EE",x"1E",x"BF",x"D0",x"F1",x"60",x"A9",x"00",x"8D",x"1C",x"BF",x"8D",x"1D",x"BF",x"A9",x"F3",x"8D",x"1E",x"BF",x"60",x"AD",x"80",x"D6",x"29",x"03",x"F0",x"13",x"EE",x"1C",x"BF",x"D0",x"0C",x"EE",x"1D",x"BF",x"D0",x"07",x"EE",x"1E",x"BF",x"D0",x"02",x"A9",x"00",x"18",x"60",x"38",x"60",x"A9",x"01",x"1C",x"30",x"D0",x"A9",x"81",x"8D",x"80",x"D6",x"38",x"60",x"48",x"A9",x"82",x"8D",x"80",x"D6",x"68",x"38",x"60",x"AD",x"80",x"D6",x"29",x"01",x"D0",x"32",x"4C",x"F3",x"A0",x"A2",x"A5",x"A0",x"AF",x"20",x"2B",x"A9",x"A2",x"F0",x"A0",x"00",x"A3",x"00",x"1B",x"D0",x"FD",x"C8",x"D0",x"FA",x"E8",x"D0",x"F7",x"A9",x"02",x"8D",x"80",x"D6",x"20",x"94",x"A0",x"20",x"A2",x"A0",x"B0",x"04",x"D0",x"F9",x"F0",x"02",x"38",x"60",x"20",x"6A",x"A0",x"4C",x"F3",x"A0",x"A9",x"07",x"8D",x"FB",x"BC",x"18",x"60",x"EE",x"81",x"D6",x"D0",x"0D",x"EE",x"82",x"D6",x"D0",x"08",x"EE",x"83",x"D6",x"D0",x"03",x"EE",x"84",x"D6",x"60",x"A9",x"01",x"8D",x"81",x"D0",x"A9",x"80",x"0C",x"86",x"D0",x"AD",x"84",x"D0",x"09",x"80",x"8D",x"7C",x"D6",x"20",x"63",x"A1",x"AD",x"85",x"D0",x"09",x"80",x"8D",x"7C",x"D6",x"20",x"63",x"A1",x"AD",x"86",x"D0",x"09",x"80",x"8D",x"7C",x"D6",x"20",x"63",x"A1",x"A9",x"21",x"8D",x"7C",x"D6",x"AD",x"86",x"D0",x"30",x"FB",x"A9",x"35",x"8D",x"AF",x"D6",x"8D",x"7F",x"D6",x"A2",x"40",x"CA",x"D0",x"FD",x"60",x"A9",x"01",x"8D",x"81",x"D0",x"A9",x"40",x"0C",x"86",x"D0",x"AD",x"84",x"D0",x"09",x"80",x"8D",x"7C",x"D6",x"20",x"63",x"A1",x"AD",x"85",x"D0",x"09",x"80",x"8D",x"7C",x"D6",x"20",x"63",x"A1",x"AD",x"86",x"D0",x"09",x"80",x"8D",x"7C",x"D6",x"20",x"63",x"A1",x"A9",x"5C",x"8D",x"7C",x"D6",x"AD",x"86",x"D0",x"29",x"C0",x"D0",x"F9",x"A9",x"16",x"8D",x"AF",x"D6",x"8D",x"7F",x"D6",x"A2",x"00",x"8A",x"20",x"69",x"A2",x"E8",x"D0",x"FA",x"A9",x"FF",x"A2",x"FE",x"20",x"84",x"A2",x"A2",x"DE",x"20",x"84",x"A2",x"A9",x"FF",x"A2",x"1E",x"20",x"84",x"A2",x"A2",x"3E",x"20",x"84",x"A2",x"20",x"55",x"A2",x"A9",x"0C",x"AA",x"A9",x"FF",x"20",x"84",x"A2",x"8A",x"18",x"69",x"20",x"90",x"F4",x"A9",x"BE",x"A2",x"C0",x"20",x"7C",x"A2",x"A2",x"D0",x"20",x"7C",x"A2",x"A2",x"F0",x"20",x"7C",x"A2",x"A2",x"E0",x"20",x"7C",x"A2",x"A2",x"00",x"20",x"7C",x"A2",x"A2",x"10",x"20",x"7C",x"A2",x"A2",x"20",x"20",x"7C",x"A2",x"A2",x"30",x"20",x"7C",x"A2",x"60",x"A2",x"C0",x"20",x"84",x"A2",x"A2",x"D0",x"20",x"84",x"A2",x"A2",x"E2",x"20",x"84",x"A2",x"A2",x"F2",x"20",x"84",x"A2",x"A2",x"00",x"20",x"84",x"A2",x"A2",x"10",x"20",x"84",x"A2",x"A2",x"22",x"20",x"84",x"A2",x"A2",x"32",x"4C",x"84",x"A2",x"A2",x"C2",x"20",x"84",x"A2",x"A2",x"D2",x"20",x"84",x"A2",x"A2",x"E0",x"20",x"84",x"A2",x"A2",x"F0",x"20",x"84",x"A2",x"A2",x"02",x"20",x"84",x"A2",x"A2",x"12",x"20",x"84",x"A2",x"A2",x"20",x"20",x"84",x"A2",x"A2",x"30",x"4C",x"84",x"A2",x"A9",x"BE",x"20",x"05",x"A2",x"A9",x"40",x"4C",x"2D",x"A2",x"A9",x"40",x"20",x"05",x"A2",x"A9",x"BE",x"4C",x"2D",x"A2",x"8E",x"F4",x"D6",x"8E",x"F4",x"D6",x"8E",x"F4",x"D6",x"8E",x"F4",x"D6",x"8E",x"F4",x"D6",x"8D",x"F5",x"D6",x"60",x"20",x"69",x"A2",x"E8",x"20",x"69",x"A2",x"E8",x"20",x"69",x"A2",x"E8",x"4C",x"69",x"A2",x"A9",x"00",x"8D",x"10",x"BF",x"A9",x"70",x"8D",x"11",x"BF",x"A9",x"FD",x"8D",x"12",x"BF",x"A9",x"0F",x"8D",x"13",x"BF",x"AD",x"29",x"D6",x"C9",x"03",x"F0",x"0A",x"AD",x"29",x"D6",x"29",x"E0",x"C9",x"20",x"F0",x"2B",x"60",x"A9",x"71",x"8D",x"11",x"BF",x"A9",x"00",x"8D",x"20",x"D0",x"A0",x"00",x"B9",x"2B",x"A3",x"C9",x"FF",x"D0",x"03",x"A3",x"00",x"60",x"4B",x"C8",x"B9",x"2B",x"A3",x"C8",x"EA",x"92",x"10",x"EE",x"20",x"D0",x"EA",x"D2",x"10",x"D0",x"F5",x"4C",x"BC",x"A2",x"A9",x"01",x"8D",x"F0",x"D6",x"A9",x"00",x"8D",x"20",x"D0",x"A0",x"00",x"B9",x"09",x"A3",x"C9",x"FF",x"D0",x"08",x"A3",x"00",x"A9",x"FF",x"8D",x"F0",x"D6",x"60",x"4B",x"C8",x"B9",x"09",x"A3",x"C8",x"EA",x"92",x"10",x"EE",x"20",x"D0",x"EA",x"D2",x"10",x"D0",x"F5",x"4C",x"E6",x"A2",x"16",x"40",x"17",x"00",x"12",x"BF",x"13",x"20",x"35",x"FF",x"36",x"FF",x"30",x"20",x"31",x"00",x"32",x"02",x"33",x"00",x"34",x"10",x"37",x"80",x"38",x"0C",x"39",x"99",x"35",x"60",x"36",x"60",x"FF",x"FF",x"E1",x"FF",x"E2",x"FF",x"DC",x"20",x"DD",x"00",x"DE",x"02",x"DF",x"00",x"E0",x"10",x"E3",x"80",x"E4",x"0C",x"E5",x"99",x"E1",x"20",x"E2",x"20",x"FF",x"FF",x"78",x"D8",x"03",x"A9",x"6B",x"8D",x"7D",x"D6",x"A9",x"02",x"0C",x"FB",x"D7",x"A9",x"3F",x"8D",x"FD",x"D7",x"20",x"A8",x"A1",x"A9",x"01",x"8D",x"FE",x"D6",x"A9",x"00",x"8D",x"1D",x"D6",x"8D",x"66",x"D0",x"8D",x"FD",x"BC",x"8D",x"1A",x"D0",x"A9",x"7F",x"8D",x"7F",x"D0",x"8D",x"0D",x"DC",x"8D",x"0D",x"DD",x"AD",x"06",x"D6",x"A9",x"40",x"8D",x"31",x"D0",x"A9",x"C5",x"0C",x"54",x"D0",x"20",x"8B",x"A2",x"A9",x"00",x"8D",x"15",x"D0",x"8D",x"63",x"D0",x"8D",x"55",x"D0",x"8D",x"6B",x"D0",x"8D",x"57",x"D0",x"A9",x"F0",x"AA",x"1C",x"49",x"D0",x"8A",x"1C",x"4B",x"D0",x"8A",x"1C",x"4D",x"D0",x"8A",x"1C",x"4F",x"D0",x"A9",x"80",x"8D",x"89",x"D6",x"20",x"CB",x"A7",x"20",x"81",x"A8",x"20",x"31",x"A8",x"60",x"78",x"A9",x"BF",x"5B",x"A0",x"BE",x"2B",x"A2",x"FF",x"9A",x"A2",x"00",x"A9",x"00",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"20",x"45",x"A3",x"20",x"34",x"A6",x"A2",x"85",x"A0",x"AE",x"20",x"2B",x"A9",x"A2",x"F7",x"A0",x"B2",x"20",x"2B",x"A9",x"A2",x"D6",x"A0",x"B2",x"20",x"2B",x"A9",x"2C",x"CB",x"A9",x"2C",x"34",x"12",x"AD",x"07",x"A4",x"C9",x"4C",x"F0",x"0A",x"A2",x"A5",x"A0",x"AE",x"20",x"2B",x"A9",x"4C",x"07",x"A4",x"A2",x"CB",x"A0",x"AE",x"20",x"2B",x"A9",x"2C",x"51",x"A4",x"20",x"CB",x"AB",x"A9",x"1A",x"8D",x"80",x"CF",x"A9",x"A4",x"8D",x"81",x"CF",x"4C",x"B3",x"AC",x"A9",x"BF",x"5B",x"A0",x"BE",x"2B",x"A2",x"FF",x"9A",x"A9",x"FF",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"01",x"0C",x"30",x"D0",x"A9",x"A9",x"8D",x"01",x"D7",x"A9",x"10",x"8D",x"05",x"D7",x"A9",x"01",x"1C",x"30",x"D0",x"A9",x"AD",x"8D",x"01",x"D7",x"A9",x"36",x"8D",x"05",x"D7",x"20",x"CB",x"A7",x"4C",x"51",x"A4",x"AD",x"10",x"D6",x"C9",x"09",x"F0",x"07",x"AD",x"11",x"D6",x"29",x"20",x"F0",x"0D",x"A2",x"48",x"A0",x"AE",x"20",x"2B",x"A9",x"EE",x"20",x"D0",x"4C",x"69",x"A4",x"20",x"81",x"A0",x"20",x"59",x"AB",x"A2",x"FF",x"20",x"2F",x"AB",x"90",x"06",x"CA",x"D0",x"F8",x"4C",x"89",x"A4",x"C9",x"1B",x"D0",x"06",x"EE",x"20",x"D0",x"4C",x"83",x"A4",x"20",x"08",x"9F",x"A2",x"2E",x"A0",x"AF",x"20",x"2B",x"A9",x"A9",x"C1",x"8D",x"80",x"D6",x"A9",x"00",x"8D",x"80",x"D6",x"A9",x"01",x"8D",x"80",x"D6",x"A2",x"03",x"20",x"81",x"A0",x"AD",x"80",x"D6",x"29",x"03",x"D0",x"0C",x"DA",x"A2",x"9F",x"A0",x"B2",x"20",x"2B",x"A9",x"FA",x"4C",x"E7",x"A4",x"CA",x"D0",x"E7",x"A9",x"C0",x"8D",x"80",x"D6",x"A2",x"8B",x"A0",x"B2",x"20",x"2B",x"A9",x"A9",x"00",x"8D",x"80",x"D6",x"A9",x"01",x"8D",x"80",x"D6",x"20",x"81",x"A0",x"AD",x"80",x"D6",x"29",x"03",x"F0",x"0A",x"A2",x"B7",x"A0",x"AF",x"20",x"2B",x"A9",x"4C",x"CB",x"A9",x"20",x"F2",x"9F",x"B0",x"1B",x"20",x"2F",x"AB",x"B0",x"07",x"C9",x"20",x"D0",x"03",x"4C",x"D6",x"AB",x"A2",x"6F",x"A0",x"AE",x"20",x"2B",x"A9",x"A9",x"81",x"0C",x"80",x"D6",x"4C",x"E7",x"A4",x"20",x"6A",x"93",x"20",x"21",x"90",x"A2",x"3C",x"A0",x"B0",x"20",x"2B",x"A9",x"A0",x"00",x"AB",x"01",x"BC",x"20",x"A4",x"A9",x"A0",x"00",x"AB",x"02",x"BC",x"20",x"A4",x"A9",x"AD",x"01",x"BC",x"D0",x"03",x"4C",x"D6",x"AB",x"20",x"CE",x"A5",x"20",x"8E",x"A6",x"A2",x"38",x"A0",x"B3",x"20",x"9C",x"99",x"20",x"99",x"98",x"B0",x"0F",x"A2",x"46",x"A0",x"B2",x"20",x"2B",x"A9",x"A0",x"00",x"AB",x"FB",x"BC",x"20",x"A4",x"A9",x"20",x"E5",x"A8",x"AD",x"7E",x"D6",x"10",x"0A",x"A2",x"0C",x"A0",x"B2",x"20",x"2B",x"A9",x"4C",x"E9",x"A5",x"A9",x"00",x"85",x"18",x"A9",x"40",x"85",x"19",x"A9",x"00",x"85",x"1A",x"A9",x"00",x"85",x"1B",x"A2",x"2D",x"A0",x"B3",x"20",x"9C",x"99",x"20",x"99",x"98",x"90",x"6E",x"A0",x"00",x"AB",x"13",x"00",x"20",x"A4",x"A9",x"AB",x"12",x"00",x"20",x"A4",x"A9",x"AB",x"11",x"00",x"20",x"A4",x"A9",x"AB",x"10",x"00",x"20",x"A4",x"A9",x"A2",x"00",x"BD",x"A3",x"A5",x"9D",x"00",x"30",x"E8",x"D0",x"F7",x"4C",x"00",x"30",x"A9",x"FF",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"A5",x"8D",x"01",x"D7",x"A9",x"BD",x"8D",x"05",x"D7",x"8D",x"7E",x"D6",x"4C",x"00",x"81",x"0A",x"80",x"00",x"81",x"FF",x"00",x"00",x"00",x"40",x"00",x"40",x"00",x"00",x"80",x"0F",x"00",x"00",x"AE",x"02",x"BC",x"20",x"D0",x"92",x"B0",x"11",x"A2",x"6B",x"A0",x"B2",x"20",x"2B",x"A9",x"A0",x"00",x"AB",x"FB",x"BC",x"20",x"A4",x"A9",x"18",x"60",x"38",x"60",x"AD",x"59",x"D6",x"29",x"01",x"D0",x"05",x"A9",x"00",x"8D",x"8B",x"D6",x"20",x"CE",x"A5",x"A9",x"50",x"8D",x"58",x"D0",x"AD",x"A1",x"D6",x"29",x"01",x"D0",x"1B",x"A2",x"1C",x"A0",x"B3",x"20",x"9C",x"99",x"20",x"DE",x"93",x"90",x"12",x"20",x"84",x"93",x"20",x"CE",x"99",x"90",x"0A",x"A2",x"4A",x"A0",x"B1",x"20",x"2B",x"A9",x"4C",x"E9",x"A6",x"A2",x"2B",x"A0",x"B1",x"20",x"2B",x"A9",x"A0",x"00",x"AB",x"FB",x"BC",x"20",x"A4",x"A9",x"4C",x"E9",x"A6",x"20",x"8E",x"A6",x"20",x"BE",x"A0",x"A9",x"00",x"A2",x"03",x"9D",x"81",x"D6",x"CA",x"10",x"FA",x"A9",x"53",x"8D",x"80",x"D6",x"CA",x"D0",x"FD",x"AD",x"71",x"DE",x"C9",x"01",x"F0",x"03",x"4C",x"CA",x"A0",x"A9",x"80",x"8D",x"82",x"D6",x"A9",x"7F",x"8D",x"83",x"D6",x"A9",x"00",x"8D",x"81",x"D6",x"8D",x"84",x"D6",x"20",x"BE",x"A0",x"A9",x"53",x"8D",x"80",x"D6",x"3A",x"10",x"FD",x"EE",x"82",x"D6",x"A2",x"00",x"A3",x"00",x"BD",x"00",x"DE",x"EA",x"92",x"18",x"1B",x"E8",x"D0",x"F6",x"E6",x"19",x"D0",x"E3",x"20",x"CA",x"A0",x"4C",x"E5",x"A8",x"A9",x"00",x"85",x"18",x"A9",x"7D",x"85",x"19",x"A9",x"05",x"85",x"1A",x"A9",x"00",x"85",x"1B",x"60",x"A2",x"04",x"A0",x"B3",x"20",x"9C",x"99",x"A9",x"00",x"85",x"18",x"A9",x"E0",x"85",x"19",x"A9",x"F7",x"85",x"1A",x"A9",x"0F",x"85",x"1B",x"4C",x"99",x"98",x"A2",x"10",x"A0",x"B3",x"20",x"9C",x"99",x"A9",x"00",x"85",x"18",x"85",x"19",x"85",x"1B",x"A9",x"02",x"85",x"1A",x"4C",x"99",x"98",x"A2",x"F8",x"A0",x"B2",x"20",x"9C",x"99",x"A9",x"00",x"85",x"18",x"A9",x"C0",x"85",x"19",x"A9",x"FD",x"85",x"1A",x"A9",x"0F",x"85",x"1B",x"4C",x"99",x"98",x"20",x"9F",x"A6",x"B0",x"03",x"4C",x"F8",x"A6",x"A2",x"09",x"A0",x"AF",x"20",x"2B",x"A9",x"20",x"B9",x"A6",x"B0",x"21",x"A2",x"0B",x"BD",x"10",x"B3",x"9D",x"C2",x"B1",x"CA",x"D0",x"F7",x"A2",x"AF",x"A0",x"B1",x"20",x"2B",x"A9",x"20",x"81",x"A0",x"20",x"81",x"A0",x"20",x"81",x"A0",x"20",x"81",x"A0",x"4C",x"B1",x"A7",x"AE",x"F9",x"BC",x"BD",x"C5",x"BC",x"8D",x"25",x"BF",x"BD",x"C6",x"BC",x"8D",x"26",x"BF",x"AD",x"26",x"BF",x"C9",x"00",x"D0",x"03",x"4C",x"9D",x"A7",x"C9",x"01",x"F0",x"F9",x"C9",x"02",x"D0",x"05",x"AD",x"25",x"BF",x"F0",x"03",x"4C",x"90",x"A7",x"20",x"09",x"85",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"00",x"A9",x"A7",x"8D",x"01",x"D7",x"A9",x"61",x"8D",x"05",x"D7",x"4C",x"70",x"A7",x"0A",x"81",x"FF",x"00",x"00",x"00",x"10",x"00",x"D0",x"02",x"00",x"E0",x"07",x"00",x"00",x"A2",x"1C",x"A0",x"AF",x"20",x"2B",x"A9",x"A2",x"EF",x"A0",x"AE",x"20",x"2B",x"A9",x"20",x"CF",x"A6",x"B0",x"07",x"A2",x"F1",x"A0",x"B1",x"20",x"2B",x"A9",x"20",x"39",x"AB",x"4C",x"CB",x"A9",x"A2",x"B8",x"A0",x"B0",x"20",x"2B",x"A9",x"20",x"81",x"A0",x"4C",x"BA",x"A3",x"A2",x"D8",x"A0",x"B0",x"20",x"2B",x"A9",x"20",x"81",x"A0",x"4C",x"BA",x"A3",x"A2",x"80",x"A0",x"B0",x"20",x"2B",x"A9",x"A2",x"8A",x"A0",x"AF",x"20",x"2B",x"A9",x"20",x"81",x"A0",x"4C",x"BA",x"A3",x"A2",x"D6",x"A0",x"AF",x"20",x"2B",x"A9",x"20",x"81",x"A0",x"4C",x"BA",x"A3",x"A9",x"40",x"8D",x"30",x"D0",x"AD",x"31",x"D0",x"29",x"40",x"8D",x"31",x"D0",x"A9",x"00",x"8D",x"20",x"D0",x"8D",x"21",x"D0",x"8D",x"11",x"D7",x"A9",x"80",x"8D",x"6F",x"D0",x"A9",x"80",x"1C",x"66",x"D0",x"A9",x"00",x"8D",x"6A",x"D0",x"8D",x"6B",x"D0",x"8D",x"78",x"D0",x"8D",x"5F",x"D0",x"A9",x"78",x"8D",x"5A",x"D0",x"A9",x"C0",x"8D",x"5D",x"D0",x"A9",x"50",x"8D",x"5C",x"D0",x"A9",x"FF",x"8D",x"01",x"DD",x"8D",x"00",x"DD",x"A9",x"14",x"8D",x"18",x"D0",x"A9",x"1B",x"8D",x"11",x"D0",x"A9",x"C8",x"8D",x"16",x"D0",x"A9",x"E5",x"8D",x"54",x"D0",x"A9",x"50",x"8D",x"58",x"D0",x"A9",x"00",x"8D",x"59",x"D0",x"60",x"A9",x"04",x"0C",x"30",x"D0",x"20",x"E5",x"A8",x"A2",x"0F",x"BD",x"51",x"A8",x"9D",x"00",x"D1",x"BD",x"61",x"A8",x"9D",x"00",x"D2",x"BD",x"71",x"A8",x"9D",x"00",x"D3",x"CA",x"10",x"EB",x"60",x"00",x"FF",x"BA",x"66",x"BB",x"55",x"D1",x"AE",x"9B",x"87",x"DD",x"B5",x"B8",x"0B",x"AA",x"8B",x"00",x"FF",x"13",x"AD",x"F3",x"EC",x"E0",x"5F",x"47",x"37",x"39",x"B5",x"B8",x"4F",x"D9",x"8B",x"00",x"FF",x"62",x"FF",x"8B",x"85",x"79",x"C7",x"81",x"00",x"78",x"B5",x"B8",x"CA",x"FE",x"8B",x"A9",x"01",x"0C",x"30",x"D0",x"A9",x"20",x"8D",x"00",x"04",x"8D",x"02",x"04",x"A9",x"00",x"8D",x"01",x"04",x"8D",x"03",x"04",x"A9",x"FF",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"A9",x"8D",x"01",x"D7",x"A9",x"10",x"8D",x"05",x"D7",x"A9",x"01",x"1C",x"30",x"D0",x"A9",x"08",x"8D",x"20",x"BF",x"A0",x"00",x"A9",x"00",x"99",x"00",x"04",x"1A",x"C8",x"C8",x"D0",x"F8",x"99",x"00",x"05",x"1A",x"C8",x"C8",x"D0",x"F8",x"99",x"00",x"06",x"1A",x"C8",x"C8",x"C0",x"80",x"D0",x"F6",x"A2",x"00",x"A9",x"16",x"9D",x"01",x"04",x"1A",x"9D",x"81",x"05",x"3A",x"9D",x"01",x"05",x"E8",x"E8",x"D0",x"F1",x"A9",x"FF",x"8D",x"70",x"D0",x"A9",x"A8",x"8D",x"01",x"D7",x"A9",x"0F",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"FF",x"8D",x"05",x"D7",x"60",x"0A",x"80",x"00",x"81",x"FF",x"00",x"00",x"00",x"03",x"00",x"7D",x"05",x"00",x"31",x"0D",x"00",x"00",x"0A",x"00",x"04",x"CC",x"07",x"00",x"04",x"00",x"04",x"04",x"00",x"00",x"00",x"81",x"FF",x"00",x"03",x"D0",x"07",x"01",x"00",x"00",x"00",x"00",x"08",x"00",x"00",x"86",x"0C",x"84",x"0D",x"A9",x"00",x"85",x"0E",x"A9",x"04",x"85",x"0F",x"AE",x"20",x"BF",x"D0",x"02",x"A2",x"08",x"E0",x"19",x"D0",x"08",x"20",x"46",x"AD",x"A2",x"18",x"8E",x"20",x"BF",x"E0",x"00",x"F0",x"10",x"18",x"A5",x"0E",x"69",x"50",x"85",x"0E",x"A5",x"0F",x"69",x"00",x"85",x"0F",x"CA",x"D0",x"EC",x"A0",x"00",x"A9",x"20",x"91",x"0E",x"C8",x"A9",x"00",x"91",x"0E",x"C8",x"C0",x"50",x"D0",x"F2",x"DB",x"A0",x"00",x"A3",x"00",x"B1",x"0C",x"F0",x"13",x"C9",x"40",x"90",x"02",x"29",x"1F",x"92",x"0E",x"1B",x"48",x"A9",x"00",x"92",x"0E",x"68",x"C8",x"1B",x"D0",x"E9",x"EE",x"20",x"BF",x"FB",x"60",x"86",x"0C",x"84",x"0D",x"A9",x"04",x"8D",x"0E",x"BF",x"A9",x"05",x"8D",x"0F",x"BF",x"20",x"6E",x"A9",x"CE",x"20",x"BF",x"60",x"6B",x"4A",x"4A",x"4A",x"4A",x"20",x"AF",x"A9",x"6B",x"29",x"0F",x"AA",x"B1",x"0E",x"C9",x"24",x"F0",x"07",x"C8",x"C8",x"C0",x"50",x"90",x"F4",x"60",x"8A",x"09",x"30",x"C9",x"3A",x"90",x"02",x"E9",x"39",x"91",x"0E",x"C8",x"C8",x"60",x"A9",x"4C",x"8D",x"D6",x"AB",x"A9",x"4C",x"8D",x"07",x"A4",x"AD",x"9D",x"D6",x"29",x"04",x"F0",x"14",x"A2",x"88",x"A0",x"B1",x"20",x"2B",x"A9",x"AD",x"10",x"D6",x"C9",x"03",x"F0",x"06",x"EE",x"20",x"D0",x"4C",x"E3",x"A9",x"8D",x"10",x"D6",x"AD",x"11",x"D6",x"29",x"04",x"F0",x"0E",x"A2",x"63",x"A0",x"B1",x"20",x"2B",x"A9",x"AD",x"11",x"D6",x"29",x"04",x"D0",x"F9",x"A9",x"82",x"8D",x"80",x"D6",x"A2",x"00",x"8A",x"9D",x"00",x"08",x"E8",x"D0",x"FA",x"A9",x"28",x"8D",x"58",x"D0",x"A9",x"00",x"8D",x"59",x"D0",x"A9",x"04",x"0C",x"7D",x"D6",x"20",x"48",x"9E",x"20",x"BD",x"9E",x"20",x"E1",x"9E",x"20",x"5D",x"AA",x"20",x"37",x"AA",x"8D",x"7F",x"D6",x"A3",x"00",x"A9",x"00",x"8D",x"10",x"BF",x"8D",x"11",x"BF",x"A9",x"01",x"8D",x"12",x"BF",x"A9",x"07",x"8D",x"13",x"BF",x"A9",x"20",x"EA",x"92",x"10",x"A0",x"00",x"1B",x"D0",x"FD",x"C8",x"D0",x"FA",x"6B",x"EA",x"92",x"10",x"60",x"AD",x"7E",x"D6",x"29",x"60",x"C9",x"40",x"F0",x"01",x"60",x"AD",x"FC",x"FF",x"8D",x"48",x"D6",x"AD",x"FD",x"FF",x"8D",x"49",x"D6",x"A9",x"AA",x"8D",x"01",x"D7",x"A9",x"0F",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"30",x"A2",x"94",x"8D",x"A0",x"AA",x"8E",x"05",x"D7",x"18",x"69",x"40",x"C9",x"30",x"D0",x"F3",x"60",x"80",x"70",x"81",x"00",x"00",x"00",x"00",x"10",x"00",x"F0",x"01",x"00",x"30",x"00",x"00",x"00",x"8E",x"CE",x"AA",x"8C",x"CF",x"AA",x"9C",x"D0",x"AA",x"8D",x"C7",x"AA",x"A9",x"AA",x"8D",x"01",x"D7",x"A9",x"0F",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"C5",x"8D",x"05",x"D7",x"60",x"0A",x"80",x"FF",x"81",x"FF",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"BC",x"0F",x"00",x"00",x"8D",x"0B",x"AB",x"8E",x"0E",x"AB",x"8C",x"0F",x"AB",x"9C",x"10",x"AB",x"6B",x"4A",x"4A",x"4A",x"4A",x"8D",x"06",x"AB",x"A9",x"01",x"8D",x"03",x"D7",x"A9",x"AB",x"8D",x"01",x"D7",x"A9",x"0F",x"8D",x"02",x"D7",x"A9",x"FF",x"8D",x"04",x"D7",x"A9",x"04",x"8D",x"05",x"D7",x"60",x"0A",x"81",x"00",x"00",x"03",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"0F",x"00",x"00",x"A9",x"00",x"A2",x"0F",x"A0",x"00",x"A3",x"3F",x"5C",x"AA",x"A0",x"00",x"A3",x"3F",x"5C",x"EA",x"60",x"AD",x"10",x"D6",x"C9",x"00",x"F0",x"02",x"18",x"60",x"38",x"60",x"20",x"24",x"AB",x"B0",x"F9",x"8D",x"10",x"D6",x"18",x"60",x"AD",x"11",x"D6",x"C9",x"20",x"F0",x"0C",x"C9",x"03",x"F0",x"05",x"29",x"10",x"D0",x"01",x"60",x"4C",x"D6",x"AB",x"AD",x"07",x"A4",x"C9",x"4C",x"F0",x"03",x"4C",x"0A",x"A4",x"4C",x"5F",x"A4",x"20",x"39",x"AB",x"A2",x"01",x"AD",x"29",x"D6",x"29",x"40",x"F0",x"02",x"A2",x"FF",x"20",x"2F",x"AB",x"90",x"06",x"CA",x"D0",x"F8",x"4C",x"7A",x"AB",x"C9",x"30",x"90",x"04",x"C9",x"39",x"90",x"02",x"A9",x"20",x"A2",x"06",x"C9",x"20",x"F0",x"04",x"9D",x"10",x"B3",x"E8",x"A9",x"2E",x"9D",x"10",x"B3",x"E8",x"A9",x"52",x"9D",x"10",x"B3",x"E8",x"A9",x"4F",x"9D",x"10",x"B3",x"E8",x"A9",x"4D",x"9D",x"10",x"B3",x"E8",x"A9",x"00",x"9D",x"10",x"B3",x"60",x"78",x"40",x"AD",x"42",x"D6",x"30",x"0E",x"C9",x"7F",x"F0",x"0A",x"8D",x"07",x"BF",x"A9",x"00",x"8D",x"06",x"BF",x"38",x"60",x"A9",x"10",x"4C",x"B1",x"92",x"A2",x"20",x"A0",x"AE",x"20",x"2B",x"A9",x"EE",x"20",x"D0",x"4C",x"C8",x"AB",x"A9",x"02",x"8D",x"1A",x"D6",x"A9",x"80",x"8D",x"6F",x"D0",x"60",x"2C",x"BE",x"AB",x"20",x"CB",x"AB",x"A2",x"D6",x"A0",x"B2",x"20",x"2B",x"A9",x"A2",x"07",x"A0",x"AE",x"20",x"2B",x"A9",x"A9",x"30",x"8D",x"08",x"BF",x"20",x"EB",x"AD",x"20",x"B3",x"AD",x"90",x"30",x"A0",x"27",x"A9",x"20",x"99",x"7A",x"AD",x"88",x"C0",x"02",x"D0",x"F8",x"C8",x"EE",x"08",x"BF",x"AD",x"08",x"BF",x"8D",x"7A",x"AD",x"A3",x"04",x"EA",x"B2",x"10",x"99",x"7A",x"AD",x"F0",x"04",x"C8",x"1B",x"80",x"F4",x"A2",x"7A",x"A0",x"AD",x"20",x"2B",x"A9",x"20",x"A2",x"AD",x"80",x"CB",x"20",x"2F",x"AB",x"C9",x"FF",x"F0",x"F9",x"C9",x"31",x"90",x"F5",x"C9",x"39",x"B0",x"F1",x"29",x"0F",x"AA",x"CA",x"20",x"EB",x"AD",x"20",x"B3",x"AD",x"90",x"E5",x"CA",x"30",x"05",x"20",x"A2",x"AD",x"80",x"F3",x"EE",x"21",x"D0",x"A3",x"24",x"EA",x"B2",x"10",x"8D",x"70",x"AD",x"1B",x"EA",x"B2",x"10",x"8D",x"71",x"AD",x"A5",x"10",x"18",x"69",x"2C",x"8D",x"72",x"AD",x"A5",x"11",x"69",x"00",x"8D",x"73",x"AD",x"20",x"D4",x"AC",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"AD",x"8D",x"01",x"D7",x"A9",x"69",x"8D",x"05",x"D7",x"A9",x"05",x"1C",x"54",x"D0",x"A9",x"28",x"8D",x"58",x"D0",x"A9",x"00",x"8D",x"59",x"D0",x"A9",x"25",x"8D",x"18",x"D0",x"A3",x"26",x"EA",x"B2",x"10",x"8D",x"48",x"D6",x"1B",x"EA",x"B2",x"10",x"8D",x"49",x"D6",x"20",x"48",x"9E",x"A9",x"3F",x"8D",x"50",x"D6",x"A9",x"36",x"8D",x"51",x"D6",x"8D",x"7F",x"D6",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"AD",x"8D",x"01",x"D7",x"A9",x"19",x"8D",x"05",x"D7",x"A9",x"00",x"5B",x"A0",x"01",x"2B",x"20",x"D4",x"AC",x"20",x"E5",x"A8",x"4C",x"0D",x"08",x"A9",x"37",x"8D",x"01",x"00",x"A9",x"97",x"1C",x"54",x"D0",x"A9",x"00",x"AA",x"A8",x"A3",x"3F",x"5C",x"EA",x"A9",x"00",x"A2",x"0F",x"5C",x"EA",x"A9",x"04",x"8D",x"88",x"02",x"AD",x"F9",x"FF",x"C9",x"FF",x"F0",x"03",x"22",x"F8",x"FF",x"A9",x"00",x"85",x"D8",x"85",x"0F",x"AD",x"7D",x"D6",x"29",x"7F",x"8D",x"7D",x"D6",x"A9",x"40",x"8D",x"20",x"04",x"A9",x"20",x"8D",x"18",x"03",x"A9",x"04",x"8D",x"19",x"03",x"60",x"0A",x"80",x"00",x"81",x"00",x"00",x"04",x"00",x"08",x"00",x"04",x"00",x"00",x"90",x"00",x"00",x"00",x"00",x"00",x"FF",x"77",x"00",x"00",x"05",x"FF",x"07",x"00",x"00",x"00",x"80",x"00",x"81",x"00",x"00",x"00",x"00",x"08",x"00",x"90",x"00",x"00",x"04",x"00",x"00",x"00",x"A9",x"FF",x"8D",x"02",x"D7",x"8D",x"04",x"D7",x"A9",x"AD",x"8D",x"01",x"D7",x"A9",x"59",x"8D",x"05",x"D7",x"60",x"80",x"00",x"81",x"00",x"00",x"00",x"00",x"05",x"D0",x"06",x"00",x"80",x"06",x"00",x"00",x"00",x"0A",x"80",x"FF",x"81",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"08",x"FF",x"07",x"00",x"00",x"00",x"31",x"2E",x"20",x"33",x"32",x"20",x"43",x"48",x"41",x"52",x"41",x"43",x"54",x"45",x"52",x"53",x"20",x"4F",x"46",x"20",x"55",x"54",x"49",x"4C",x"49",x"54",x"59",x"20",x"4E",x"41",x"4D",x"45",x"2E",x"2E",x"2E",x"20",x"20",x"20",x"20",x"00",x"A3",x"2A",x"EA",x"B2",x"10",x"DA",x"AA",x"1B",x"EA",x"B2",x"10",x"85",x"11",x"86",x"10",x"FA",x"60",x"A3",x"00",x"EA",x"B2",x"10",x"C9",x"4D",x"D0",x"2D",x"1B",x"EA",x"B2",x"10",x"C9",x"36",x"D0",x"25",x"1B",x"EA",x"B2",x"10",x"C9",x"35",x"D0",x"1D",x"1B",x"EA",x"B2",x"10",x"C9",x"55",x"D0",x"15",x"A3",x"28",x"EA",x"B2",x"10",x"CD",x"10",x"BF",x"D0",x"0B",x"1B",x"EA",x"B2",x"10",x"CD",x"11",x"BF",x"D0",x"02",x"38",x"60",x"18",x"60",x"A9",x"50",x"85",x"10",x"A9",x"08",x"85",x"11",x"A9",x"F8",x"85",x"12",x"A9",x"0F",x"85",x"13",x"60",x"AE",x"7C",x"D6",x"D0",x"FB",x"8D",x"7C",x"D6",x"8D",x"7F",x"D6",x"53",x"45",x"4C",x"45",x"43",x"54",x"20",x"55",x"54",x"49",x"4C",x"49",x"54",x"59",x"20",x"54",x"4F",x"20",x"4C",x"41",x"55",x"4E",x"43",x"48",x"00",x"48",x"4F",x"4C",x"44",x"20",x"41",x"4C",x"54",x"20",x"2B",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"43",x"59",x"43",x"4C",x"45",x"20",x"46",x"4F",x"52",x"20",x"55",x"54",x"49",x"4C",x"49",x"54",x"59",x"20",x"4D",x"45",x"4E",x"55",x"00",x"48",x"4F",x"4C",x"44",x"20",x"4E",x"4F",x"20",x"53",x"43",x"52",x"4F",x"4C",x"4C",x"20",x"2B",x"20",x"50",x"4F",x"57",x"45",x"52",x"20",x"43",x"59",x"43",x"4C",x"45",x"20",x"46",x"4F",x"52",x"20",x"46",x"4C",x"41",x"53",x"48",x"00",x"52",x"45",x"2D",x"54",x"52",x"59",x"49",x"4E",x"47",x"20",x"54",x"4F",x"20",x"52",x"45",x"41",x"44",x"20",x"4D",x"42",x"52",x"00",x"4D",x"45",x"47",x"41",x"36",x"35",x"20",x"4D",x"45",x"47",x"41",x"4F",x"53",x"20",x"48",x"59",x"50",x"45",x"52",x"56",x"49",x"53",x"4F",x"52",x"20",x"56",x"30",x"30",x"2E",x"31",x"37",x"00",x"4E",x"4F",x"20",x"53",x"43",x"52",x"4F",x"4C",x"4C",x"3D",x"46",x"4C",x"41",x"53",x"48",x"2C",x"20",x"41",x"4C",x"54",x"3D",x"55",x"54",x"49",x"4C",x"53",x"2C",x"20",x"43",x"54",x"52",x"4C",x"3D",x"48",x"4F",x"4C",x"44",x"00",x"50",x"4F",x"57",x"45",x"52",x"20",x"4F",x"46",x"46",x"2F",x"4F",x"4E",x"20",x"46",x"4F",x"52",x"20",x"46",x"4C",x"41",x"53",x"48",x"20",x"4F",x"52",x"20",x"55",x"54",x"49",x"4C",x"20",x"4D",x"45",x"4E",x"55",x"00",x"52",x"4F",x"4D",x"20",x"43",x"48",x"45",x"43",x"4B",x"53",x"55",x"4D",x"20",x"4F",x"4B",x"20",x"2D",x"20",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"00",x"4C",x"4F",x"41",x"44",x"45",x"44",x"20",x"43",x"48",x"41",x"52",x"52",x"4F",x"4D",x"2E",x"4D",x"36",x"35",x"00",x"4C",x"4F",x"41",x"44",x"45",x"44",x"20",x"4D",x"45",x"47",x"41",x"36",x"35",x"2E",x"52",x"4F",x"4D",x"00",x"4C",x"4F",x"4F",x"4B",x"49",x"4E",x"47",x"20",x"46",x"4F",x"52",x"20",x"53",x"44",x"48",x"43",x"20",x"43",x"41",x"52",x"44",x"20",x"3E",x"3D",x"34",x"47",x"42",x"2E",x"2E",x"2E",x"00",x"53",x"44",x"20",x"43",x"41",x"52",x"44",x"20",x"49",x"53",x"20",x"4E",x"4F",x"54",x"20",x"53",x"44",x"48",x"43",x"2E",x"20",x"4D",x"55",x"53",x"54",x"20",x"42",x"45",x"20",x"53",x"44",x"48",x"43",x"2E",x"00",x"46",x"4F",x"55",x"4E",x"44",x"20",x"41",x"4E",x"44",x"20",x"52",x"45",x"53",x"45",x"54",x"20",x"53",x"44",x"48",x"43",x"20",x"43",x"41",x"52",x"44",x"00",x"45",x"52",x"52",x"4F",x"52",x"20",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53",x"44",x"20",x"43",x"41",x"52",x"44",x"00",x"52",x"45",x"2D",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"00",x"4E",x"4F",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"2C",x"20",x"54",x"52",x"59",x"49",x"4E",x"47",x"20",x"42",x"55",x"49",x"4C",x"54",x"2D",x"49",x"4E",x"20",x"52",x"4F",x"4D",x"00",x"42",x"41",x"44",x"20",x"4D",x"42",x"52",x"20",x"4F",x"52",x"20",x"44",x"4F",x"53",x"20",x"42",x"4F",x"4F",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"2E",x"00",x"52",x"45",x"41",x"44",x"20",x"50",x"41",x"52",x"54",x"49",x"54",x"49",x"4F",x"4E",x"20",x"54",x"41",x"42",x"4C",x"45",x"20",x"46",x"52",x"4F",x"4D",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"00",x"46",x"4F",x"55",x"4E",x"44",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"2E",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"43",x"4C",x"55",x"53",x"54",x"45",x"52",x"20",x"3D",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"44",x"49",x"53",x"4B",x"2D",x"43",x"4F",x"55",x"4E",x"54",x"3D",x"24",x"24",x"2C",x"20",x"44",x"45",x"46",x"41",x"55",x"4C",x"54",x"2D",x"44",x"49",x"53",x"4B",x"3D",x"24",x"24",x"00",x"4C",x"4F",x"4F",x"4B",x"49",x"4E",x"47",x"20",x"46",x"4F",x"52",x"20",x"24",x"24",x"20",x"42",x"59",x"54",x"45",x"53",x"2C",x"20",x"49",x"20",x"53",x"45",x"45",x"20",x"24",x"24",x"20",x"42",x"59",x"54",x"45",x"53",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"4F",x"50",x"45",x"4E",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"20",x"46",x"4F",x"52",x"20",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"00",x"52",x"45",x"41",x"44",x"49",x"4E",x"47",x"20",x"52",x"4F",x"4D",x"20",x"46",x"49",x"4C",x"45",x"2E",x"2E",x"2E",x"00",x"52",x"4F",x"4D",x"20",x"54",x"4F",x"4F",x"20",x"4C",x"4F",x"4E",x"47",x"3A",x"20",x"28",x"52",x"45",x"41",x"44",x"20",x"24",x"24",x"24",x"24",x"20",x"50",x"41",x"47",x"45",x"53",x"29",x"00",x"52",x"4F",x"4D",x"20",x"54",x"4F",x"4F",x"20",x"53",x"48",x"4F",x"52",x"54",x"3A",x"20",x"28",x"52",x"45",x"41",x"44",x"20",x"24",x"24",x"24",x"24",x"20",x"50",x"41",x"47",x"45",x"53",x"29",x"00",x"43",x"55",x"52",x"52",x"45",x"4E",x"54",x"20",x"43",x"4C",x"55",x"53",x"54",x"45",x"52",x"3D",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"43",x"55",x"52",x"52",x"45",x"4E",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"3D",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"43",x"41",x"4E",x"4E",x"4F",x"54",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"20",x"44",x"38",x"31",x"20",x"2D",x"20",x"28",x"45",x"52",x"52",x"4E",x"4F",x"3A",x"20",x"24",x"24",x"29",x"00",x"44",x"38",x"31",x"20",x"53",x"55",x"43",x"43",x"45",x"53",x"53",x"46",x"55",x"4C",x"4C",x"59",x"20",x"4D",x"4F",x"55",x"4E",x"54",x"45",x"44",x"00",x"52",x"45",x"4C",x"45",x"41",x"53",x"45",x"20",x"43",x"4F",x"4E",x"54",x"52",x"4F",x"4C",x"20",x"54",x"4F",x"20",x"43",x"4F",x"4E",x"54",x"49",x"4E",x"55",x"45",x"20",x"42",x"4F",x"4F",x"54",x"49",x"4E",x"47",x"2E",x"00",x"53",x"57",x"33",x"20",x"4F",x"46",x"46",x"20",x"4F",x"52",x"20",x"50",x"52",x"45",x"53",x"53",x"20",x"52",x"55",x"4E",x"2F",x"53",x"54",x"4F",x"50",x"20",x"54",x"4F",x"20",x"43",x"4F",x"4E",x"54",x"49",x"4E",x"55",x"45",x"2E",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"46",x"49",x"4E",x"44",x"20",x"52",x"4F",x"4D",x"20",x"4D",x"45",x"47",x"41",x"36",x"35",x"58",x"58",x"52",x"4F",x"4D",x"00",x"4C",x"4F",x"41",x"44",x"49",x"4E",x"47",x"20",x"48",x"49",x"43",x"4B",x"55",x"50",x"2E",x"4D",x"36",x"35",x"20",x"49",x"4E",x"54",x"4F",x"20",x"48",x"59",x"50",x"45",x"52",x"56",x"49",x"53",x"4F",x"52",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"4C",x"4F",x"41",x"44",x"20",x"31",x"35",x"34",x"31",x"52",x"4F",x"4D",x"2E",x"4D",x"36",x"35",x"00",x"52",x"55",x"4E",x"4E",x"49",x"4E",x"47",x"20",x"48",x"49",x"43",x"4B",x"45",x"44",x"20",x"48",x"59",x"50",x"45",x"52",x"56",x"49",x"53",x"4F",x"52",x"00",x"4C",x"4F",x"4F",x"4B",x"49",x"4E",x"47",x"20",x"46",x"4F",x"52",x"20",x"4E",x"45",x"58",x"54",x"20",x"53",x"45",x"43",x"54",x"4F",x"52",x"20",x"4F",x"46",x"20",x"46",x"49",x"4C",x"45",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"4C",x"4F",x"41",x"44",x"20",x"42",x"41",x"4E",x"4E",x"45",x"52",x"2E",x"4D",x"36",x"35",x"20",x"28",x"45",x"52",x"52",x"4E",x"4F",x"3A",x"24",x"24",x"29",x"00",x"43",x"4F",x"55",x"4C",x"44",x"20",x"4E",x"4F",x"54",x"20",x"43",x"48",x"44",x"49",x"52",x"20",x"54",x"4F",x"20",x"2F",x"20",x"28",x"45",x"52",x"52",x"4E",x"4F",x"3A",x"24",x"24",x"29",x"00",x"54",x"52",x"59",x"49",x"4E",x"47",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"42",x"55",x"53",x"20",x"30",x"00",x"55",x"53",x"49",x"4E",x"47",x"20",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"42",x"55",x"53",x"20",x"31",x"00",x"44",x"4D",x"41",x"47",x"49",x"43",x"20",x"52",x"45",x"56",x"20",x"41",x"20",x"4D",x"4F",x"44",x"45",x"00",x"44",x"4D",x"41",x"47",x"49",x"43",x"20",x"52",x"45",x"56",x"20",x"42",x"20",x"4D",x"4F",x"44",x"45",x"00",x"47",x"49",x"54",x"3A",x"20",x"6D",x"61",x"73",x"74",x"65",x"72",x"2C",x"32",x"30",x"32",x"33",x"31",x"30",x"30",x"35",x"2E",x"31",x"32",x"2C",x"66",x"39",x"33",x"38",x"35",x"37",x"30",x"7E",x"00",x"00",x"31",x"35",x"34",x"31",x"52",x"4F",x"4D",x"2E",x"4D",x"36",x"35",x"00",x"43",x"48",x"41",x"52",x"52",x"4F",x"4D",x"2E",x"4D",x"36",x"35",x"00",x"4D",x"45",x"47",x"41",x"36",x"35",x"2E",x"52",x"4F",x"4D",x"00",x"00",x"4D",x"45",x"47",x"41",x"36",x"35",x"2E",x"44",x"38",x"31",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"48",x"49",x"43",x"4B",x"55",x"50",x"2E",x"4D",x"36",x"35",x"00",x"42",x"41",x"4E",x"4E",x"45",x"52",x"2E",x"4D",x"36",x"35",x"00",x"46",x"52",x"45",x"45",x"5A",x"45",x"52",x"2E",x"4D",x"36",x"35",x"00",x"4E",x"54",x"53",x"43",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"56",x"65",x"6E",x"65",x"7A",x"75",x"61",x"6C",x"65",x"6E",x"20",x"63",x"61",x"73",x"61",x"62",x"61",x"20",x"6D",x"65",x"6C",x"6F",x"6E",x"20",x"70",x"72",x"6F",x"64",x"75",x"63",x"74",x"69",x"6F",x"6E",x"20",x"73",x"74",x"61",x"74",x"69",x"73",x"74",x"69",x"63",x"73",x"20",x"28",x"32",x"30",x"31",x"32",x"2D",x"32",x"30",x"31",x"35",x"29",x"2E",x"74",x"78",x"74",x"20",x"20",x"00",x"00",x"46",x"49",x"4C",x"45",x"4E",x"41",x"4D",x"45",x"2E",x"45",x"58",x"54",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"56",x"65",x"6E",x"65",x"7A",x"75",x"61",x"6C",x"65",x"6E",x"20",x"63",x"61",x"73",x"61",x"62",x"61",x"20",x"6D",x"65",x"6C",x"6F",x"6E",x"20",x"70",x"72",x"6F",x"64",x"75",x"63",x"74",x"69",x"6F",x"6E",x"20",x"73",x"74",x"61",x"74",x"69",x"73",x"74",x"69",x"63",x"73",x"20",x"28",x"32",x"30",x"30",x"37",x"2D",x"32",x"30",x"31",x"31",x"29",x"2E",x"74",x"78",x"74",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"4F",x"50",x"45",x"52",x"41",x"54",x"49",x"4E",x"47",x"20",x"53",x"59",x"53",x"54",x"45",x"4D",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");

begin

--process for read and write operation.
  PROCESS(Clk,cs,ram,address,address_i)
  BEGIN
    if(rising_edge(Clk)) then 
      if cs='1' then
        if(we='1') then
          ram(to_integer(unsigned(address_i))) <= data_i;
        end if;
      end if;
      data_o <= ram(to_integer(unsigned(address)));
    end if;
--    if cs='1' then
--      data_o <= ram(to_integer(unsigned(address)));
--    else
--      data_o <= "ZZZZZZZZ";
--    end if;
  END PROCESS;

end Behavioral;
