--------------------------------------------------------------------------------
--                              Compressor_23_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          X1 : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3 is
signal X :  std_logic_vector(4 downto 0);
begin
   X <=X1 & X0 ;
   with X select R <= 
      "000" when "00000", 
      "001" when "00001", 
      "001" when "00010", 
      "010" when "00011", 
      "001" when "00100", 
      "010" when "00101", 
      "010" when "00110", 
      "011" when "00111", 
      "010" when "01000", 
      "011" when "01001", 
      "011" when "01010", 
      "100" when "01011", 
      "011" when "01100", 
      "100" when "01101", 
      "100" when "01110", 
      "101" when "01111", 
      "010" when "10000", 
      "011" when "10001", 
      "011" when "10010", 
      "100" when "10011", 
      "011" when "10100", 
      "100" when "10101", 
      "100" when "10110", 
      "101" when "10111", 
      "100" when "11000", 
      "101" when "11001", 
      "101" when "11010", 
      "110" when "11011", 
      "101" when "11100", 
      "110" when "11101", 
      "110" when "11110", 
      "111" when "11111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                             LZOC_46_F400_uid4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_46_F400_uid4 is
   port ( clk, rst : in std_logic;
          I : in  std_logic_vector(45 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of LZOC_46_F400_uid4 is
signal sozb, sozb_d1, sozb_d2, sozb_d3 :  std_logic;
signal level6, level6_d1 :  std_logic_vector(63 downto 0);
signal digit6, digit6_d1, digit6_d2, digit6_d3 :  std_logic;
signal level5 :  std_logic_vector(31 downto 0);
signal digit5, digit5_d1, digit5_d2 :  std_logic;
signal level4, level4_d1 :  std_logic_vector(15 downto 0);
signal digit4, digit4_d1 :  std_logic;
signal level3 :  std_logic_vector(7 downto 0);
signal digit3, digit3_d1 :  std_logic;
signal level2, level2_d1 :  std_logic_vector(3 downto 0);
signal digit2 :  std_logic;
signal level1 :  std_logic_vector(1 downto 0);
signal digit1 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            sozb_d3 <=  sozb_d2;
            level6_d1 <=  level6;
            digit6_d1 <=  digit6;
            digit6_d2 <=  digit6_d1;
            digit6_d3 <=  digit6_d2;
            digit5_d1 <=  digit5;
            digit5_d2 <=  digit5_d1;
            level4_d1 <=  level4;
            digit4_d1 <=  digit4;
            digit3_d1 <=  digit3;
            level2_d1 <=  level2;
         end if;
      end process;
   sozb <= OZB;
   level6<= I& (17 downto 0 => not(sozb));
   digit6<= '1' when level6(63 downto 32) = (63 downto 32 => sozb) else '0';
   ----------------Synchro barrier, entering cycle 1----------------
   level5<= level6_d1(31 downto 0) when digit6_d1='1' else level6_d1(63 downto 32);
   digit5<= '1' when level5(31 downto 16) = (31 downto 16 => sozb_d1) else '0';
   level4<= level5(15 downto 0) when digit5='1' else level5(31 downto 16);
   ----------------Synchro barrier, entering cycle 2----------------
   digit4<= '1' when level4_d1(15 downto 8) = (15 downto 8 => sozb_d2) else '0';
   level3<= level4_d1(7 downto 0) when digit4='1' else level4_d1(15 downto 8);
   digit3<= '1' when level3(7 downto 4) = (7 downto 4 => sozb_d2) else '0';
   level2<= level3(3 downto 0) when digit3='1' else level3(7 downto 4);
   ----------------Synchro barrier, entering cycle 3----------------
   digit2<= '1' when level2_d1(3 downto 2) = (3 downto 2 => sozb_d3) else '0';
   level1<= level2_d1(1 downto 0) when digit2='1' else level2_d1(3 downto 2);
   digit1<= '1' when level1(1 downto 1) = (1 downto 1 => sozb_d3) else '0';
   O <= digit6_d3 & digit5_d2 & digit4_d1 & digit3_d1 & digit2 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                     LeftShifter_24_by_max_24_F400_uid8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_24_by_max_24_F400_uid8 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(23 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(47 downto 0)   );
end entity;

architecture arch of LeftShifter_24_by_max_24_F400_uid8 is
signal level0 :  std_logic_vector(23 downto 0);
signal ps, ps_d1 :  std_logic_vector(4 downto 0);
signal level1 :  std_logic_vector(24 downto 0);
signal level2, level2_d1 :  std_logic_vector(26 downto 0);
signal level3 :  std_logic_vector(30 downto 0);
signal level4 :  std_logic_vector(38 downto 0);
signal level5 :  std_logic_vector(54 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level2_d1 <=  level2;
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   ----------------Synchro barrier, entering cycle 1----------------
   level3<= level2_d1 & (3 downto 0 => '0') when ps_d1(2)= '1' else     (3 downto 0 => '0') & level2_d1;
   level4<= level3 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps_d1(4)= '1' else     (15 downto 0 => '0') & level4;
   R <= level5(47 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        InvTable_0_10_11_F400_uid12
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity InvTable_0_10_11_F400_uid12 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(10 downto 0)   );
end entity;

architecture arch of InvTable_0_10_11_F400_uid12 is
signal TableOut, TableOut_d1 :  std_logic_vector(10 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            TableOut_d1 <=  TableOut;
         end if;
      end process;
  with X select TableOut <= 
   "10000000000" when "0000000000",
   "10000000000" when "0000000001",
   "01111111111" when "0000000010",
   "01111111110" when "0000000011",
   "01111111101" when "0000000100",
   "01111111100" when "0000000101",
   "01111111011" when "0000000110",
   "01111111010" when "0000000111",
   "01111111001" when "0000001000",
   "01111111000" when "0000001001",
   "01111110111" when "0000001010",
   "01111110110" when "0000001011",
   "01111110101" when "0000001100",
   "01111110100" when "0000001101",
   "01111110011" when "0000001110",
   "01111110010" when "0000001111",
   "01111110001" when "0000010000",
   "01111110000" when "0000010001",
   "01111101111" when "0000010010",
   "01111101110" when "0000010011",
   "01111101101" when "0000010100",
   "01111101100" when "0000010101",
   "01111101011" when "0000010110",
   "01111101010" when "0000010111",
   "01111101001" when "0000011000",
   "01111101000" when "0000011001",
   "01111100111" when "0000011010",
   "01111100110" when "0000011011",
   "01111100101" when "0000011100",
   "01111100100" when "0000011101",
   "01111100011" when "0000011110",
   "01111100010" when "0000011111",
   "01111100001" when "0000100000",
   "01111100001" when "0000100001",
   "01111100000" when "0000100010",
   "01111011111" when "0000100011",
   "01111011110" when "0000100100",
   "01111011101" when "0000100101",
   "01111011100" when "0000100110",
   "01111011011" when "0000100111",
   "01111011010" when "0000101000",
   "01111011001" when "0000101001",
   "01111011000" when "0000101010",
   "01111010111" when "0000101011",
   "01111010110" when "0000101100",
   "01111010101" when "0000101101",
   "01111010100" when "0000101110",
   "01111010100" when "0000101111",
   "01111010011" when "0000110000",
   "01111010010" when "0000110001",
   "01111010001" when "0000110010",
   "01111010000" when "0000110011",
   "01111001111" when "0000110100",
   "01111001110" when "0000110101",
   "01111001101" when "0000110110",
   "01111001100" when "0000110111",
   "01111001011" when "0000111000",
   "01111001011" when "0000111001",
   "01111001010" when "0000111010",
   "01111001001" when "0000111011",
   "01111001000" when "0000111100",
   "01111000111" when "0000111101",
   "01111000110" when "0000111110",
   "01111000101" when "0000111111",
   "01111000100" when "0001000000",
   "01111000011" when "0001000001",
   "01111000010" when "0001000010",
   "01111000010" when "0001000011",
   "01111000001" when "0001000100",
   "01111000000" when "0001000101",
   "01110111111" when "0001000110",
   "01110111110" when "0001000111",
   "01110111101" when "0001001000",
   "01110111100" when "0001001001",
   "01110111011" when "0001001010",
   "01110111011" when "0001001011",
   "01110111010" when "0001001100",
   "01110111001" when "0001001101",
   "01110111000" when "0001001110",
   "01110110111" when "0001001111",
   "01110110110" when "0001010000",
   "01110110101" when "0001010001",
   "01110110101" when "0001010010",
   "01110110100" when "0001010011",
   "01110110011" when "0001010100",
   "01110110010" when "0001010101",
   "01110110001" when "0001010110",
   "01110110000" when "0001010111",
   "01110101111" when "0001011000",
   "01110101111" when "0001011001",
   "01110101110" when "0001011010",
   "01110101101" when "0001011011",
   "01110101100" when "0001011100",
   "01110101011" when "0001011101",
   "01110101010" when "0001011110",
   "01110101010" when "0001011111",
   "01110101001" when "0001100000",
   "01110101000" when "0001100001",
   "01110100111" when "0001100010",
   "01110100110" when "0001100011",
   "01110100101" when "0001100100",
   "01110100101" when "0001100101",
   "01110100100" when "0001100110",
   "01110100011" when "0001100111",
   "01110100010" when "0001101000",
   "01110100001" when "0001101001",
   "01110100000" when "0001101010",
   "01110100000" when "0001101011",
   "01110011111" when "0001101100",
   "01110011110" when "0001101101",
   "01110011101" when "0001101110",
   "01110011100" when "0001101111",
   "01110011100" when "0001110000",
   "01110011011" when "0001110001",
   "01110011010" when "0001110010",
   "01110011001" when "0001110011",
   "01110011000" when "0001110100",
   "01110010111" when "0001110101",
   "01110010111" when "0001110110",
   "01110010110" when "0001110111",
   "01110010101" when "0001111000",
   "01110010100" when "0001111001",
   "01110010011" when "0001111010",
   "01110010011" when "0001111011",
   "01110010010" when "0001111100",
   "01110010001" when "0001111101",
   "01110010000" when "0001111110",
   "01110010000" when "0001111111",
   "01110001111" when "0010000000",
   "01110001110" when "0010000001",
   "01110001101" when "0010000010",
   "01110001100" when "0010000011",
   "01110001100" when "0010000100",
   "01110001011" when "0010000101",
   "01110001010" when "0010000110",
   "01110001001" when "0010000111",
   "01110001000" when "0010001000",
   "01110001000" when "0010001001",
   "01110000111" when "0010001010",
   "01110000110" when "0010001011",
   "01110000101" when "0010001100",
   "01110000101" when "0010001101",
   "01110000100" when "0010001110",
   "01110000011" when "0010001111",
   "01110000010" when "0010010000",
   "01110000001" when "0010010001",
   "01110000001" when "0010010010",
   "01110000000" when "0010010011",
   "01101111111" when "0010010100",
   "01101111110" when "0010010101",
   "01101111110" when "0010010110",
   "01101111101" when "0010010111",
   "01101111100" when "0010011000",
   "01101111011" when "0010011001",
   "01101111011" when "0010011010",
   "01101111010" when "0010011011",
   "01101111001" when "0010011100",
   "01101111000" when "0010011101",
   "01101111000" when "0010011110",
   "01101110111" when "0010011111",
   "01101110110" when "0010100000",
   "01101110101" when "0010100001",
   "01101110101" when "0010100010",
   "01101110100" when "0010100011",
   "01101110011" when "0010100100",
   "01101110010" when "0010100101",
   "01101110010" when "0010100110",
   "01101110001" when "0010100111",
   "01101110000" when "0010101000",
   "01101101111" when "0010101001",
   "01101101111" when "0010101010",
   "01101101110" when "0010101011",
   "01101101101" when "0010101100",
   "01101101101" when "0010101101",
   "01101101100" when "0010101110",
   "01101101011" when "0010101111",
   "01101101010" when "0010110000",
   "01101101010" when "0010110001",
   "01101101001" when "0010110010",
   "01101101000" when "0010110011",
   "01101100111" when "0010110100",
   "01101100111" when "0010110101",
   "01101100110" when "0010110110",
   "01101100101" when "0010110111",
   "01101100101" when "0010111000",
   "01101100100" when "0010111001",
   "01101100011" when "0010111010",
   "01101100010" when "0010111011",
   "01101100010" when "0010111100",
   "01101100001" when "0010111101",
   "01101100000" when "0010111110",
   "01101100000" when "0010111111",
   "01101011111" when "0011000000",
   "01101011110" when "0011000001",
   "01101011101" when "0011000010",
   "01101011101" when "0011000011",
   "01101011100" when "0011000100",
   "01101011011" when "0011000101",
   "01101011011" when "0011000110",
   "01101011010" when "0011000111",
   "01101011001" when "0011001000",
   "01101011000" when "0011001001",
   "01101011000" when "0011001010",
   "01101010111" when "0011001011",
   "01101010110" when "0011001100",
   "01101010110" when "0011001101",
   "01101010101" when "0011001110",
   "01101010100" when "0011001111",
   "01101010100" when "0011010000",
   "01101010011" when "0011010001",
   "01101010010" when "0011010010",
   "01101010010" when "0011010011",
   "01101010001" when "0011010100",
   "01101010000" when "0011010101",
   "01101001111" when "0011010110",
   "01101001111" when "0011010111",
   "01101001110" when "0011011000",
   "01101001101" when "0011011001",
   "01101001101" when "0011011010",
   "01101001100" when "0011011011",
   "01101001011" when "0011011100",
   "01101001011" when "0011011101",
   "01101001010" when "0011011110",
   "01101001001" when "0011011111",
   "01101001001" when "0011100000",
   "01101001000" when "0011100001",
   "01101000111" when "0011100010",
   "01101000111" when "0011100011",
   "01101000110" when "0011100100",
   "01101000101" when "0011100101",
   "01101000101" when "0011100110",
   "01101000100" when "0011100111",
   "01101000011" when "0011101000",
   "01101000011" when "0011101001",
   "01101000010" when "0011101010",
   "01101000001" when "0011101011",
   "01101000001" when "0011101100",
   "01101000000" when "0011101101",
   "01100111111" when "0011101110",
   "01100111111" when "0011101111",
   "01100111110" when "0011110000",
   "01100111101" when "0011110001",
   "01100111101" when "0011110010",
   "01100111100" when "0011110011",
   "01100111011" when "0011110100",
   "01100111011" when "0011110101",
   "01100111010" when "0011110110",
   "01100111010" when "0011110111",
   "01100111001" when "0011111000",
   "01100111000" when "0011111001",
   "01100111000" when "0011111010",
   "01100110111" when "0011111011",
   "01100110110" when "0011111100",
   "01100110110" when "0011111101",
   "01100110101" when "0011111110",
   "01100110100" when "0011111111",
   "01100110100" when "0100000000",
   "01100110011" when "0100000001",
   "01100110010" when "0100000010",
   "01100110010" when "0100000011",
   "01100110001" when "0100000100",
   "01100110001" when "0100000101",
   "01100110000" when "0100000110",
   "01100101111" when "0100000111",
   "01100101111" when "0100001000",
   "01100101110" when "0100001001",
   "01100101101" when "0100001010",
   "01100101101" when "0100001011",
   "01100101100" when "0100001100",
   "01100101011" when "0100001101",
   "01100101011" when "0100001110",
   "01100101010" when "0100001111",
   "01100101010" when "0100010000",
   "01100101001" when "0100010001",
   "01100101000" when "0100010010",
   "01100101000" when "0100010011",
   "01100100111" when "0100010100",
   "01100100110" when "0100010101",
   "01100100110" when "0100010110",
   "01100100101" when "0100010111",
   "01100100101" when "0100011000",
   "01100100100" when "0100011001",
   "01100100011" when "0100011010",
   "01100100011" when "0100011011",
   "01100100010" when "0100011100",
   "01100100010" when "0100011101",
   "01100100001" when "0100011110",
   "01100100000" when "0100011111",
   "01100100000" when "0100100000",
   "01100011111" when "0100100001",
   "01100011111" when "0100100010",
   "01100011110" when "0100100011",
   "01100011101" when "0100100100",
   "01100011101" when "0100100101",
   "01100011100" when "0100100110",
   "01100011011" when "0100100111",
   "01100011011" when "0100101000",
   "01100011010" when "0100101001",
   "01100011010" when "0100101010",
   "01100011001" when "0100101011",
   "01100011000" when "0100101100",
   "01100011000" when "0100101101",
   "01100010111" when "0100101110",
   "01100010111" when "0100101111",
   "01100010110" when "0100110000",
   "01100010101" when "0100110001",
   "01100010101" when "0100110010",
   "01100010100" when "0100110011",
   "01100010100" when "0100110100",
   "01100010011" when "0100110101",
   "01100010011" when "0100110110",
   "01100010010" when "0100110111",
   "01100010001" when "0100111000",
   "01100010001" when "0100111001",
   "01100010000" when "0100111010",
   "01100010000" when "0100111011",
   "01100001111" when "0100111100",
   "01100001110" when "0100111101",
   "01100001110" when "0100111110",
   "01100001101" when "0100111111",
   "01100001101" when "0101000000",
   "01100001100" when "0101000001",
   "01100001100" when "0101000010",
   "01100001011" when "0101000011",
   "01100001010" when "0101000100",
   "01100001010" when "0101000101",
   "01100001001" when "0101000110",
   "01100001001" when "0101000111",
   "01100001000" when "0101001000",
   "01100001000" when "0101001001",
   "01100000111" when "0101001010",
   "01100000110" when "0101001011",
   "01100000110" when "0101001100",
   "01100000101" when "0101001101",
   "01100000101" when "0101001110",
   "01100000100" when "0101001111",
   "01100000100" when "0101010000",
   "01100000011" when "0101010001",
   "01100000010" when "0101010010",
   "01100000010" when "0101010011",
   "01100000001" when "0101010100",
   "01100000001" when "0101010101",
   "01100000000" when "0101010110",
   "01100000000" when "0101010111",
   "01011111111" when "0101011000",
   "01011111110" when "0101011001",
   "01011111110" when "0101011010",
   "01011111101" when "0101011011",
   "01011111101" when "0101011100",
   "01011111100" when "0101011101",
   "01011111100" when "0101011110",
   "01011111011" when "0101011111",
   "01011111011" when "0101100000",
   "01011111010" when "0101100001",
   "01011111001" when "0101100010",
   "01011111001" when "0101100011",
   "01011111000" when "0101100100",
   "01011111000" when "0101100101",
   "01011110111" when "0101100110",
   "01011110111" when "0101100111",
   "01011110110" when "0101101000",
   "01011110110" when "0101101001",
   "01011110101" when "0101101010",
   "01011110101" when "0101101011",
   "01011110100" when "0101101100",
   "01011110011" when "0101101101",
   "01011110011" when "0101101110",
   "01011110010" when "0101101111",
   "01011110010" when "0101110000",
   "01011110001" when "0101110001",
   "01011110001" when "0101110010",
   "01011110000" when "0101110011",
   "01011110000" when "0101110100",
   "01011101111" when "0101110101",
   "01011101111" when "0101110110",
   "01011101110" when "0101110111",
   "01011101101" when "0101111000",
   "01011101101" when "0101111001",
   "01011101100" when "0101111010",
   "01011101100" when "0101111011",
   "01011101011" when "0101111100",
   "01011101011" when "0101111101",
   "01011101010" when "0101111110",
   "01011101010" when "0101111111",
   "01011101001" when "0110000000",
   "01011101001" when "0110000001",
   "01011101000" when "0110000010",
   "01011101000" when "0110000011",
   "01011100111" when "0110000100",
   "01011100111" when "0110000101",
   "01011100110" when "0110000110",
   "01011100110" when "0110000111",
   "01011100101" when "0110001000",
   "01011100100" when "0110001001",
   "01011100100" when "0110001010",
   "01011100011" when "0110001011",
   "01011100011" when "0110001100",
   "01011100010" when "0110001101",
   "01011100010" when "0110001110",
   "01011100001" when "0110001111",
   "01011100001" when "0110010000",
   "01011100000" when "0110010001",
   "01011100000" when "0110010010",
   "01011011111" when "0110010011",
   "01011011111" when "0110010100",
   "01011011110" when "0110010101",
   "01011011110" when "0110010110",
   "01011011101" when "0110010111",
   "01011011101" when "0110011000",
   "01011011100" when "0110011001",
   "01011011100" when "0110011010",
   "01011011011" when "0110011011",
   "01011011011" when "0110011100",
   "01011011010" when "0110011101",
   "01011011010" when "0110011110",
   "01011011001" when "0110011111",
   "01011011001" when "0110100000",
   "01011011000" when "0110100001",
   "01011011000" when "0110100010",
   "01011010111" when "0110100011",
   "01011010111" when "0110100100",
   "01011010110" when "0110100101",
   "01011010110" when "0110100110",
   "01011010101" when "0110100111",
   "01011010101" when "0110101000",
   "01011010100" when "0110101001",
   "01011010100" when "0110101010",
   "01011010011" when "0110101011",
   "01011010011" when "0110101100",
   "01011010010" when "0110101101",
   "01011010010" when "0110101110",
   "01011010001" when "0110101111",
   "01011010001" when "0110110000",
   "01011010000" when "0110110001",
   "01011010000" when "0110110010",
   "01011001111" when "0110110011",
   "01011001111" when "0110110100",
   "01011001110" when "0110110101",
   "01011001110" when "0110110110",
   "01011001101" when "0110110111",
   "01011001101" when "0110111000",
   "01011001100" when "0110111001",
   "01011001100" when "0110111010",
   "01011001011" when "0110111011",
   "01011001011" when "0110111100",
   "01011001010" when "0110111101",
   "01011001010" when "0110111110",
   "01011001001" when "0110111111",
   "01011001001" when "0111000000",
   "01011001000" when "0111000001",
   "01011001000" when "0111000010",
   "01011000111" when "0111000011",
   "01011000111" when "0111000100",
   "01011000110" when "0111000101",
   "01011000110" when "0111000110",
   "01011000101" when "0111000111",
   "01011000101" when "0111001000",
   "01011000101" when "0111001001",
   "01011000100" when "0111001010",
   "01011000100" when "0111001011",
   "01011000011" when "0111001100",
   "01011000011" when "0111001101",
   "01011000010" when "0111001110",
   "01011000010" when "0111001111",
   "01011000001" when "0111010000",
   "01011000001" when "0111010001",
   "01011000000" when "0111010010",
   "01011000000" when "0111010011",
   "01010111111" when "0111010100",
   "01010111111" when "0111010101",
   "01010111110" when "0111010110",
   "01010111110" when "0111010111",
   "01010111101" when "0111011000",
   "01010111101" when "0111011001",
   "01010111100" when "0111011010",
   "01010111100" when "0111011011",
   "01010111100" when "0111011100",
   "01010111011" when "0111011101",
   "01010111011" when "0111011110",
   "01010111010" when "0111011111",
   "01010111010" when "0111100000",
   "01010111001" when "0111100001",
   "01010111001" when "0111100010",
   "01010111000" when "0111100011",
   "01010111000" when "0111100100",
   "01010110111" when "0111100101",
   "01010110111" when "0111100110",
   "01010110110" when "0111100111",
   "01010110110" when "0111101000",
   "01010110110" when "0111101001",
   "01010110101" when "0111101010",
   "01010110101" when "0111101011",
   "01010110100" when "0111101100",
   "01010110100" when "0111101101",
   "01010110011" when "0111101110",
   "01010110011" when "0111101111",
   "01010110010" when "0111110000",
   "01010110010" when "0111110001",
   "01010110001" when "0111110010",
   "01010110001" when "0111110011",
   "01010110001" when "0111110100",
   "01010110000" when "0111110101",
   "01010110000" when "0111110110",
   "01010101111" when "0111110111",
   "01010101111" when "0111111000",
   "01010101110" when "0111111001",
   "01010101110" when "0111111010",
   "01010101101" when "0111111011",
   "01010101101" when "0111111100",
   "01010101101" when "0111111101",
   "01010101100" when "0111111110",
   "01010101100" when "0111111111",
   "10101010110" when "1000000000",
   "10101010101" when "1000000001",
   "10101010100" when "1000000010",
   "10101010011" when "1000000011",
   "10101010010" when "1000000100",
   "10101010001" when "1000000101",
   "10101010001" when "1000000110",
   "10101010000" when "1000000111",
   "10101001111" when "1000001000",
   "10101001110" when "1000001001",
   "10101001101" when "1000001010",
   "10101001100" when "1000001011",
   "10101001011" when "1000001100",
   "10101001010" when "1000001101",
   "10101001010" when "1000001110",
   "10101001001" when "1000001111",
   "10101001000" when "1000010000",
   "10101000111" when "1000010001",
   "10101000110" when "1000010010",
   "10101000101" when "1000010011",
   "10101000100" when "1000010100",
   "10101000011" when "1000010101",
   "10101000011" when "1000010110",
   "10101000010" when "1000010111",
   "10101000001" when "1000011000",
   "10101000000" when "1000011001",
   "10100111111" when "1000011010",
   "10100111110" when "1000011011",
   "10100111101" when "1000011100",
   "10100111101" when "1000011101",
   "10100111100" when "1000011110",
   "10100111011" when "1000011111",
   "10100111010" when "1000100000",
   "10100111001" when "1000100001",
   "10100111000" when "1000100010",
   "10100110111" when "1000100011",
   "10100110111" when "1000100100",
   "10100110110" when "1000100101",
   "10100110101" when "1000100110",
   "10100110100" when "1000100111",
   "10100110011" when "1000101000",
   "10100110010" when "1000101001",
   "10100110001" when "1000101010",
   "10100110001" when "1000101011",
   "10100110000" when "1000101100",
   "10100101111" when "1000101101",
   "10100101110" when "1000101110",
   "10100101101" when "1000101111",
   "10100101100" when "1000110000",
   "10100101100" when "1000110001",
   "10100101011" when "1000110010",
   "10100101010" when "1000110011",
   "10100101001" when "1000110100",
   "10100101000" when "1000110101",
   "10100100111" when "1000110110",
   "10100100111" when "1000110111",
   "10100100110" when "1000111000",
   "10100100101" when "1000111001",
   "10100100100" when "1000111010",
   "10100100011" when "1000111011",
   "10100100011" when "1000111100",
   "10100100010" when "1000111101",
   "10100100001" when "1000111110",
   "10100100000" when "1000111111",
   "10100011111" when "1001000000",
   "10100011110" when "1001000001",
   "10100011110" when "1001000010",
   "10100011101" when "1001000011",
   "10100011100" when "1001000100",
   "10100011011" when "1001000101",
   "10100011010" when "1001000110",
   "10100011010" when "1001000111",
   "10100011001" when "1001001000",
   "10100011000" when "1001001001",
   "10100010111" when "1001001010",
   "10100010110" when "1001001011",
   "10100010101" when "1001001100",
   "10100010101" when "1001001101",
   "10100010100" when "1001001110",
   "10100010011" when "1001001111",
   "10100010010" when "1001010000",
   "10100010001" when "1001010001",
   "10100010001" when "1001010010",
   "10100010000" when "1001010011",
   "10100001111" when "1001010100",
   "10100001110" when "1001010101",
   "10100001101" when "1001010110",
   "10100001101" when "1001010111",
   "10100001100" when "1001011000",
   "10100001011" when "1001011001",
   "10100001010" when "1001011010",
   "10100001001" when "1001011011",
   "10100001001" when "1001011100",
   "10100001000" when "1001011101",
   "10100000111" when "1001011110",
   "10100000110" when "1001011111",
   "10100000110" when "1001100000",
   "10100000101" when "1001100001",
   "10100000100" when "1001100010",
   "10100000011" when "1001100011",
   "10100000010" when "1001100100",
   "10100000010" when "1001100101",
   "10100000001" when "1001100110",
   "10100000000" when "1001100111",
   "10011111111" when "1001101000",
   "10011111110" when "1001101001",
   "10011111110" when "1001101010",
   "10011111101" when "1001101011",
   "10011111100" when "1001101100",
   "10011111011" when "1001101101",
   "10011111011" when "1001101110",
   "10011111010" when "1001101111",
   "10011111001" when "1001110000",
   "10011111000" when "1001110001",
   "10011111000" when "1001110010",
   "10011110111" when "1001110011",
   "10011110110" when "1001110100",
   "10011110101" when "1001110101",
   "10011110100" when "1001110110",
   "10011110100" when "1001110111",
   "10011110011" when "1001111000",
   "10011110010" when "1001111001",
   "10011110001" when "1001111010",
   "10011110001" when "1001111011",
   "10011110000" when "1001111100",
   "10011101111" when "1001111101",
   "10011101110" when "1001111110",
   "10011101110" when "1001111111",
   "10011101101" when "1010000000",
   "10011101100" when "1010000001",
   "10011101011" when "1010000010",
   "10011101011" when "1010000011",
   "10011101010" when "1010000100",
   "10011101001" when "1010000101",
   "10011101000" when "1010000110",
   "10011101000" when "1010000111",
   "10011100111" when "1010001000",
   "10011100110" when "1010001001",
   "10011100101" when "1010001010",
   "10011100101" when "1010001011",
   "10011100100" when "1010001100",
   "10011100011" when "1010001101",
   "10011100010" when "1010001110",
   "10011100010" when "1010001111",
   "10011100001" when "1010010000",
   "10011100000" when "1010010001",
   "10011011111" when "1010010010",
   "10011011111" when "1010010011",
   "10011011110" when "1010010100",
   "10011011101" when "1010010101",
   "10011011100" when "1010010110",
   "10011011100" when "1010010111",
   "10011011011" when "1010011000",
   "10011011010" when "1010011001",
   "10011011001" when "1010011010",
   "10011011001" when "1010011011",
   "10011011000" when "1010011100",
   "10011010111" when "1010011101",
   "10011010110" when "1010011110",
   "10011010110" when "1010011111",
   "10011010101" when "1010100000",
   "10011010100" when "1010100001",
   "10011010100" when "1010100010",
   "10011010011" when "1010100011",
   "10011010010" when "1010100100",
   "10011010001" when "1010100101",
   "10011010001" when "1010100110",
   "10011010000" when "1010100111",
   "10011001111" when "1010101000",
   "10011001111" when "1010101001",
   "10011001110" when "1010101010",
   "10011001101" when "1010101011",
   "10011001100" when "1010101100",
   "10011001100" when "1010101101",
   "10011001011" when "1010101110",
   "10011001010" when "1010101111",
   "10011001001" when "1010110000",
   "10011001001" when "1010110001",
   "10011001000" when "1010110010",
   "10011000111" when "1010110011",
   "10011000111" when "1010110100",
   "10011000110" when "1010110101",
   "10011000101" when "1010110110",
   "10011000100" when "1010110111",
   "10011000100" when "1010111000",
   "10011000011" when "1010111001",
   "10011000010" when "1010111010",
   "10011000010" when "1010111011",
   "10011000001" when "1010111100",
   "10011000000" when "1010111101",
   "10011000000" when "1010111110",
   "10010111111" when "1010111111",
   "10010111110" when "1011000000",
   "10010111101" when "1011000001",
   "10010111101" when "1011000010",
   "10010111100" when "1011000011",
   "10010111011" when "1011000100",
   "10010111011" when "1011000101",
   "10010111010" when "1011000110",
   "10010111001" when "1011000111",
   "10010111001" when "1011001000",
   "10010111000" when "1011001001",
   "10010110111" when "1011001010",
   "10010110110" when "1011001011",
   "10010110110" when "1011001100",
   "10010110101" when "1011001101",
   "10010110100" when "1011001110",
   "10010110100" when "1011001111",
   "10010110011" when "1011010000",
   "10010110010" when "1011010001",
   "10010110010" when "1011010010",
   "10010110001" when "1011010011",
   "10010110000" when "1011010100",
   "10010110000" when "1011010101",
   "10010101111" when "1011010110",
   "10010101110" when "1011010111",
   "10010101110" when "1011011000",
   "10010101101" when "1011011001",
   "10010101100" when "1011011010",
   "10010101011" when "1011011011",
   "10010101011" when "1011011100",
   "10010101010" when "1011011101",
   "10010101001" when "1011011110",
   "10010101001" when "1011011111",
   "10010101000" when "1011100000",
   "10010100111" when "1011100001",
   "10010100111" when "1011100010",
   "10010100110" when "1011100011",
   "10010100101" when "1011100100",
   "10010100101" when "1011100101",
   "10010100100" when "1011100110",
   "10010100011" when "1011100111",
   "10010100011" when "1011101000",
   "10010100010" when "1011101001",
   "10010100001" when "1011101010",
   "10010100001" when "1011101011",
   "10010100000" when "1011101100",
   "10010011111" when "1011101101",
   "10010011111" when "1011101110",
   "10010011110" when "1011101111",
   "10010011101" when "1011110000",
   "10010011101" when "1011110001",
   "10010011100" when "1011110010",
   "10010011011" when "1011110011",
   "10010011011" when "1011110100",
   "10010011010" when "1011110101",
   "10010011001" when "1011110110",
   "10010011001" when "1011110111",
   "10010011000" when "1011111000",
   "10010010111" when "1011111001",
   "10010010111" when "1011111010",
   "10010010110" when "1011111011",
   "10010010101" when "1011111100",
   "10010010101" when "1011111101",
   "10010010100" when "1011111110",
   "10010010011" when "1011111111",
   "10010010011" when "1100000000",
   "10010010010" when "1100000001",
   "10010010001" when "1100000010",
   "10010010001" when "1100000011",
   "10010010000" when "1100000100",
   "10010010000" when "1100000101",
   "10010001111" when "1100000110",
   "10010001110" when "1100000111",
   "10010001110" when "1100001000",
   "10010001101" when "1100001001",
   "10010001100" when "1100001010",
   "10010001100" when "1100001011",
   "10010001011" when "1100001100",
   "10010001010" when "1100001101",
   "10010001010" when "1100001110",
   "10010001001" when "1100001111",
   "10010001000" when "1100010000",
   "10010001000" when "1100010001",
   "10010000111" when "1100010010",
   "10010000111" when "1100010011",
   "10010000110" when "1100010100",
   "10010000101" when "1100010101",
   "10010000101" when "1100010110",
   "10010000100" when "1100010111",
   "10010000011" when "1100011000",
   "10010000011" when "1100011001",
   "10010000010" when "1100011010",
   "10010000001" when "1100011011",
   "10010000001" when "1100011100",
   "10010000000" when "1100011101",
   "10010000000" when "1100011110",
   "10001111111" when "1100011111",
   "10001111110" when "1100100000",
   "10001111110" when "1100100001",
   "10001111101" when "1100100010",
   "10001111100" when "1100100011",
   "10001111100" when "1100100100",
   "10001111011" when "1100100101",
   "10001111010" when "1100100110",
   "10001111010" when "1100100111",
   "10001111001" when "1100101000",
   "10001111001" when "1100101001",
   "10001111000" when "1100101010",
   "10001110111" when "1100101011",
   "10001110111" when "1100101100",
   "10001110110" when "1100101101",
   "10001110101" when "1100101110",
   "10001110101" when "1100101111",
   "10001110100" when "1100110000",
   "10001110100" when "1100110001",
   "10001110011" when "1100110010",
   "10001110010" when "1100110011",
   "10001110010" when "1100110100",
   "10001110001" when "1100110101",
   "10001110001" when "1100110110",
   "10001110000" when "1100110111",
   "10001101111" when "1100111000",
   "10001101111" when "1100111001",
   "10001101110" when "1100111010",
   "10001101101" when "1100111011",
   "10001101101" when "1100111100",
   "10001101100" when "1100111101",
   "10001101100" when "1100111110",
   "10001101011" when "1100111111",
   "10001101010" when "1101000000",
   "10001101010" when "1101000001",
   "10001101001" when "1101000010",
   "10001101001" when "1101000011",
   "10001101000" when "1101000100",
   "10001100111" when "1101000101",
   "10001100111" when "1101000110",
   "10001100110" when "1101000111",
   "10001100110" when "1101001000",
   "10001100101" when "1101001001",
   "10001100100" when "1101001010",
   "10001100100" when "1101001011",
   "10001100011" when "1101001100",
   "10001100011" when "1101001101",
   "10001100010" when "1101001110",
   "10001100001" when "1101001111",
   "10001100001" when "1101010000",
   "10001100000" when "1101010001",
   "10001100000" when "1101010010",
   "10001011111" when "1101010011",
   "10001011110" when "1101010100",
   "10001011110" when "1101010101",
   "10001011101" when "1101010110",
   "10001011101" when "1101010111",
   "10001011100" when "1101011000",
   "10001011011" when "1101011001",
   "10001011011" when "1101011010",
   "10001011010" when "1101011011",
   "10001011010" when "1101011100",
   "10001011001" when "1101011101",
   "10001011000" when "1101011110",
   "10001011000" when "1101011111",
   "10001010111" when "1101100000",
   "10001010111" when "1101100001",
   "10001010110" when "1101100010",
   "10001010110" when "1101100011",
   "10001010101" when "1101100100",
   "10001010100" when "1101100101",
   "10001010100" when "1101100110",
   "10001010011" when "1101100111",
   "10001010011" when "1101101000",
   "10001010010" when "1101101001",
   "10001010001" when "1101101010",
   "10001010001" when "1101101011",
   "10001010000" when "1101101100",
   "10001010000" when "1101101101",
   "10001001111" when "1101101110",
   "10001001111" when "1101101111",
   "10001001110" when "1101110000",
   "10001001101" when "1101110001",
   "10001001101" when "1101110010",
   "10001001100" when "1101110011",
   "10001001100" when "1101110100",
   "10001001011" when "1101110101",
   "10001001010" when "1101110110",
   "10001001010" when "1101110111",
   "10001001001" when "1101111000",
   "10001001001" when "1101111001",
   "10001001000" when "1101111010",
   "10001001000" when "1101111011",
   "10001000111" when "1101111100",
   "10001000110" when "1101111101",
   "10001000110" when "1101111110",
   "10001000101" when "1101111111",
   "10001000101" when "1110000000",
   "10001000100" when "1110000001",
   "10001000100" when "1110000010",
   "10001000011" when "1110000011",
   "10001000010" when "1110000100",
   "10001000010" when "1110000101",
   "10001000001" when "1110000110",
   "10001000001" when "1110000111",
   "10001000000" when "1110001000",
   "10001000000" when "1110001001",
   "10000111111" when "1110001010",
   "10000111111" when "1110001011",
   "10000111110" when "1110001100",
   "10000111101" when "1110001101",
   "10000111101" when "1110001110",
   "10000111100" when "1110001111",
   "10000111100" when "1110010000",
   "10000111011" when "1110010001",
   "10000111011" when "1110010010",
   "10000111010" when "1110010011",
   "10000111010" when "1110010100",
   "10000111001" when "1110010101",
   "10000111000" when "1110010110",
   "10000111000" when "1110010111",
   "10000110111" when "1110011000",
   "10000110111" when "1110011001",
   "10000110110" when "1110011010",
   "10000110110" when "1110011011",
   "10000110101" when "1110011100",
   "10000110101" when "1110011101",
   "10000110100" when "1110011110",
   "10000110011" when "1110011111",
   "10000110011" when "1110100000",
   "10000110010" when "1110100001",
   "10000110010" when "1110100010",
   "10000110001" when "1110100011",
   "10000110001" when "1110100100",
   "10000110000" when "1110100101",
   "10000110000" when "1110100110",
   "10000101111" when "1110100111",
   "10000101110" when "1110101000",
   "10000101110" when "1110101001",
   "10000101101" when "1110101010",
   "10000101101" when "1110101011",
   "10000101100" when "1110101100",
   "10000101100" when "1110101101",
   "10000101011" when "1110101110",
   "10000101011" when "1110101111",
   "10000101010" when "1110110000",
   "10000101010" when "1110110001",
   "10000101001" when "1110110010",
   "10000101001" when "1110110011",
   "10000101000" when "1110110100",
   "10000100111" when "1110110101",
   "10000100111" when "1110110110",
   "10000100110" when "1110110111",
   "10000100110" when "1110111000",
   "10000100101" when "1110111001",
   "10000100101" when "1110111010",
   "10000100100" when "1110111011",
   "10000100100" when "1110111100",
   "10000100011" when "1110111101",
   "10000100011" when "1110111110",
   "10000100010" when "1110111111",
   "10000100010" when "1111000000",
   "10000100001" when "1111000001",
   "10000100000" when "1111000010",
   "10000100000" when "1111000011",
   "10000011111" when "1111000100",
   "10000011111" when "1111000101",
   "10000011110" when "1111000110",
   "10000011110" when "1111000111",
   "10000011101" when "1111001000",
   "10000011101" when "1111001001",
   "10000011100" when "1111001010",
   "10000011100" when "1111001011",
   "10000011011" when "1111001100",
   "10000011011" when "1111001101",
   "10000011010" when "1111001110",
   "10000011010" when "1111001111",
   "10000011001" when "1111010000",
   "10000011001" when "1111010001",
   "10000011000" when "1111010010",
   "10000011000" when "1111010011",
   "10000010111" when "1111010100",
   "10000010110" when "1111010101",
   "10000010110" when "1111010110",
   "10000010101" when "1111010111",
   "10000010101" when "1111011000",
   "10000010100" when "1111011001",
   "10000010100" when "1111011010",
   "10000010011" when "1111011011",
   "10000010011" when "1111011100",
   "10000010010" when "1111011101",
   "10000010010" when "1111011110",
   "10000010001" when "1111011111",
   "10000010001" when "1111100000",
   "10000010000" when "1111100001",
   "10000010000" when "1111100010",
   "10000001111" when "1111100011",
   "10000001111" when "1111100100",
   "10000001110" when "1111100101",
   "10000001110" when "1111100110",
   "10000001101" when "1111100111",
   "10000001101" when "1111101000",
   "10000001100" when "1111101001",
   "10000001100" when "1111101010",
   "10000001011" when "1111101011",
   "10000001011" when "1111101100",
   "10000001010" when "1111101101",
   "10000001010" when "1111101110",
   "10000001001" when "1111101111",
   "10000001001" when "1111110000",
   "10000001000" when "1111110001",
   "10000001000" when "1111110010",
   "10000000111" when "1111110011",
   "10000000111" when "1111110100",
   "10000000110" when "1111110101",
   "10000000110" when "1111110110",
   "10000000101" when "1111110111",
   "10000000101" when "1111111000",
   "10000000100" when "1111111001",
   "10000000100" when "1111111010",
   "10000000011" when "1111111011",
   "10000000011" when "1111111100",
   "10000000010" when "1111111101",
   "10000000010" when "1111111110",
   "10000000001" when "1111111111",
   "-----------" when others;
    Y <= TableOut_d1;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_59_f400_uid16
--                    (IntAdderAlternative_59_F400_uid20)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_59_f400_uid16 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(58 downto 0);
          Y : in  std_logic_vector(58 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(58 downto 0)   );
end entity;

architecture arch of IntAdder_59_f400_uid16 is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(17 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(16 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(17 downto 0);
signal sum_l1_idx1 :  std_logic_vector(16 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(58 downto 42)) + ( "0" & Y(58 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
   sum_l0_idx1 <= s_sum_l0_idx1(16 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(17 downto 17);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(16 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(17 downto 17);
   R <= sum_l1_idx1(16 downto 0) & sum_l0_idx0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_59_f400_uid24
--                    (IntAdderAlternative_59_F400_uid28)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_59_f400_uid24 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(58 downto 0);
          Y : in  std_logic_vector(58 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(58 downto 0)   );
end entity;

architecture arch of IntAdder_59_f400_uid24 is
signal s_sum_l0_idx0 :  std_logic_vector(33 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(26 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(32 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(25 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(26 downto 0);
signal sum_l1_idx1 :  std_logic_vector(25 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(32 downto 0)) + ( "0" & Y(32 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(58 downto 33)) + ( "0" & Y(58 downto 33));
   sum_l0_idx0 <= s_sum_l0_idx0(32 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(33 downto 33);
   sum_l0_idx1 <= s_sum_l0_idx1(25 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(26 downto 26);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(25 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(26 downto 26);
   R <= sum_l1_idx1(25 downto 0) & sum_l0_idx0_d1(32 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_50_f400_uid32
--                     (IntAdderClassical_50_F400_uid34)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_50_f400_uid32 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(49 downto 0);
          Y : in  std_logic_vector(49 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of IntAdder_50_f400_uid32 is
signal x0 :  std_logic_vector(23 downto 0);
signal y0 :  std_logic_vector(23 downto 0);
signal x1, x1_d1 :  std_logic_vector(25 downto 0);
signal y1, y1_d1 :  std_logic_vector(25 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(24 downto 0);
signal sum1 :  std_logic_vector(26 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
         end if;
      end process;
   --Classical
   x0 <= X(23 downto 0);
   y0 <= Y(23 downto 0);
   x1 <= X(49 downto 24);
   y1 <= Y(49 downto 24);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin;
   ----------------Synchro barrier, entering cycle 1----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(24);
   R <= sum1(25 downto 0) & sum0_d1(23 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_50_f400_uid40
--                     (IntAdderClassical_50_F400_uid42)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_50_f400_uid40 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(49 downto 0);
          Y : in  std_logic_vector(49 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of IntAdder_50_f400_uid40 is
signal x0 :  std_logic_vector(23 downto 0);
signal y0 :  std_logic_vector(23 downto 0);
signal x1, x1_d1 :  std_logic_vector(25 downto 0);
signal y1, y1_d1 :  std_logic_vector(25 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(24 downto 0);
signal sum1 :  std_logic_vector(26 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
         end if;
      end process;
   --Classical
   x0 <= X(23 downto 0);
   y0 <= Y(23 downto 0);
   x1 <= X(49 downto 24);
   y1 <= Y(49 downto 24);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin;
   ----------------Synchro barrier, entering cycle 1----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(24);
   R <= sum1(25 downto 0) & sum0_d1(23 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntSquarer_28_F400_uid48
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2009)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee; 
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
library work;
entity IntSquarer_28_F400_uid48 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          R : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of IntSquarer_28_F400_uid48 is
signal x0_16, x0_16_d1, x0_16_d2 :  std_logic_vector(17 downto 0);
signal x17_32, x17_32_d1, x17_32_d2, x17_32_d3 :  std_logic_vector(17 downto 0);
signal x17_32_shr, x17_32_shr_d1, x17_32_shr_d2 :  std_logic_vector(17 downto 0);
signal p0, p0_d1, p0_d2 :  std_logic_vector(35 downto 0);
signal p1_x2, p1_x2_d1 :  std_logic_vector(35 downto 0);
signal s1, s1_d1 :  std_logic_vector(35 downto 0);
signal p2, p2_d1 :  std_logic_vector(35 downto 0);
signal s2 :  std_logic_vector(35 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            x0_16_d1 <=  x0_16;
            x0_16_d2 <=  x0_16_d1;
            x17_32_d1 <=  x17_32;
            x17_32_d2 <=  x17_32_d1;
            x17_32_d3 <=  x17_32_d2;
            x17_32_shr_d1 <=  x17_32_shr;
            x17_32_shr_d2 <=  x17_32_shr_d1;
            p0_d1 <=  p0;
            p0_d2 <=  p0_d1;
            p1_x2_d1 <=  p1_x2;
            s1_d1 <=  s1;
            p2_d1 <=  p2;
         end if;
      end process;
   x0_16 <= "0" & X(16 downto 0);
   x17_32 <= "00" & "00000" & X(27 downto 17);
   x17_32_shr <= "0" & "00000" & X(27 downto 17) & "0";
   ----------------Synchro barrier, entering cycle 1----------------
   ----------------Synchro barrier, entering cycle 2----------------
   p0 <= x0_16_d2 * x0_16_d2;
   p1_x2 <= x17_32_shr_d2 * x0_16_d2;
   ----------------Synchro barrier, entering cycle 3----------------
   s1 <= p1_x2_d1 + ( "00000000000000000" & p0_d1(35 downto 17));
   p2 <= x17_32_d3 * x17_32_d3;
   ----------------Synchro barrier, entering cycle 4----------------
   s2 <= p2_d1 + ( "00000000000000000" & s1_d1(35 downto 17));
   R <= s2(21 downto 0) & s1_d1(16 downto 0) & p0_d2(16 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_50_f400_uid52
--                     (IntAdderClassical_50_F400_uid54)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_50_f400_uid52 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(49 downto 0);
          Y : in  std_logic_vector(49 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(49 downto 0)   );
end entity;

architecture arch of IntAdder_50_f400_uid52 is
signal x0 :  std_logic_vector(21 downto 0);
signal y0 :  std_logic_vector(21 downto 0);
signal x1, x1_d1 :  std_logic_vector(27 downto 0);
signal y1, y1_d1 :  std_logic_vector(27 downto 0);
signal sum0, sum0_d1 :  std_logic_vector(22 downto 0);
signal sum1 :  std_logic_vector(28 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            sum0_d1 <=  sum0;
         end if;
      end process;
   --Classical
   x0 <= X(21 downto 0);
   y0 <= Y(21 downto 0);
   x1 <= X(49 downto 22);
   y1 <= Y(49 downto 22);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin;
   ----------------Synchro barrier, entering cycle 1----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(22);
   R <= sum1(27 downto 0) & sum0_d1(21 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        LogTable_0_10_74_F400_uid60
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity LogTable_0_10_74_F400_uid60 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(73 downto 0)   );
end entity;

architecture arch of LogTable_0_10_74_F400_uid60 is
signal TableOut, TableOut_d1 :  std_logic_vector(73 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            TableOut_d1 <=  TableOut;
         end if;
      end process;
  with X select TableOut <= 
   "11111111111111101111111111111100000000000000000000000000000000000000000000" when "0000000000",
   "11111111111111101111111111111100000000000000000000000000000000000000000000" when "0000000001",
   "00000000001111110000011111111101010101011001010101100010001001001100110101" when "0000000010",
   "00000000011111110010000000000110101011101010110001000100111011110011100001" when "0000000011",
   "00000000101111110100100000100000000101000100110000101110000000110100101101" when "0000000100",
   "00000000111111111000000001010001100101011000100010110011010101111110010110" when "0000000101",
   "00000001001111111100100010100011010001111000011110001110000111000111011111" when "0000000110",
   "00000001100000000010000100011101010001011000011010110101010000001110000011" when "0000000111",
   "00000001110000001000100111000111101100001110001001111111101010101110110111" when "0000001000",
   "00000010000000010000001010101010101100010001101111001110001001010001100110" when "0000001001",
   "00000010010000011000101111001110011100111101111000111101000100100011100011" when "0000001010",
   "00000010100000100010010100111011001011010000011001011101111100011101010110" when "0000001011",
   "00000010110000101100111011111001000101101010011111111000110000010001010100" when "0000001100",
   "00000011000000111000100100010000011100010001010001010101010001000001001011" when "0000001101",
   "00000011010001000101001110001001100000101110000010001100010000111011001010" when "0000001110",
   "00000011100001010010111001101100100110001110101111100000110011000000001100" when "0000001111",
   "00000011110001100001100111000010000001100110011000100001011101110101110001" when "0000010000",
   "00000100000001110001010110010010001001001101011000010001110100100111110010" when "0000010001",
   "00000100010010000010000111100101010101000001111111011011111001011111111011" when "0000010010",
   "00000100100010010011111011000011111110101000101110001001111100011001010001" when "0000010011",
   "00000100110010100110110000110110100001001100101110001000011001011000100110" when "0000010100",
   "00000101000010111010101001000101011001100000001100110000001001110011001001" when "0000010101",
   "00000101010011001111100011111001000101111100110101011001001011001110100110" when "0000010110",
   "00000101100011100101100001011010000110100100001011110101011111100111000101" when "0000010111",
   "00000101110011111100100001110000111101000000000110110100101001101001000100" when "0000011000",
   "00000110000100010100100101000110001100100011001010101111101000101110011011" when "0000011001",
   "00000110010100101101101011100010011010001001000100011101010111101111100110" when "0000011010",
   "00000110100101000111110101001110001100010111000100001111110001111011000010" when "0000011011",
   "00000110110101100011000010010010001011011100011000111001100001000110111001" when "0000011100",
   "00000111000101111111010010110111000001010010101010111100011000110001111111" when "0000011101",
   "00000111010110011100100111000101011001011110011000000000100001001010111101" when "0000011110",
   "00000111100110111010111111000110000001001111001110010100010101110101101101" when "0000011111",
   "00000111110111011010011011000001100111100000101000010101011011001001001110" when "0000100000",
   "00000111110111011010011011000001100111100000101000010101011011001001001110" when "0000100001",
   "00001000000111111010111011000000111100111010001000100010001110000000101110" when "0000100010",
   "00001000011000011100011111001100110011101111110101010100110001011101010100" when "0000100011",
   "00001000101000111111000111101110000000000010110101000110011101010110010111" when "0000100100",
   "00001000111001100010110100101101010111100001101010011100110001111000110110" when "0000100101",
   "00001001001010000111100110010011110001101000110000011111010011010111000000" when "0000100110",
   "00001001011010101101011100101010000111100010110111010110110001101011101010" when "0000100111",
   "00001001101011010100010111111001010100001001100000110101011111010101111100" when "0000101000",
   "00001001111011111100011000001010010100000101011101001000111011010011111110" when "0000101001",
   "00001010001100100101011101100110000101101111000111110100110001100100010100" when "0000101010",
   "00001010011101001111101000010101101001001111000100110111010101111000010010" when "0000101011",
   "00001010101101111010111000100010000000011110011101110111011100100010000001" when "0000101100",
   "00001010111110100111001110010100001111000111011111011011110100101100000000" when "0000101101",
   "00001011001111010100101001110101011010100101110110101100001000001000001010" when "0000101110",
   "00001011001111010100101001110101011010100101110110101100001000001000001010" when "0000101111",
   "00001011100000000011001011001110101010000111001110111011100100000111011100" when "0000110000",
   "00001011110000110010110010101001000110101011101111011101001111001011111000" when "0000110001",
   "00001100000001100011100000001101111011000110011001100010001111101001000011" when "0000110010",
   "00001100010010010101010100000110010011111101100110100001100110101000110000" when "0000110011",
   "00001100100011001000001110011011011111101011100110001010000011101011000001" when "0000110100",
   "00001100110011111100001111010110101110011110111100111101110100011011000101" when "0000110101",
   "00001101000100110001010111000001010010011011000010111000010100110011111110" when "0000110110",
   "00001101010101100111100101100100011111011000100001111110000011010001101010" when "0000110111",
   "00001101100110011110111011001001101011000101110101010110011101001101011011" when "0000111000",
   "00001101100110011110111011001001101011000101110101010110011101001101011011" when "0000111001",
   "00001101110111010111010111111010001101000111101000010000000111100101110100" when "0000111010",
   "00001110001000010000111011111111011110111001010101001111000111110100100110" when "0000111011",
   "00001110011001001011100111100010111011101101100101100101110000110110111000" when "0000111100",
   "00001110101010000111011010101110000000101110110000110111101000101101010111" when "0000111101",
   "00001110111011000100010101101010001100111111011100100111001010011100110110" when "0000111110",
   "00001111001100000010011000100001000001011010111100001101101000111000101110" when "0000111111",
   "00001111011101000001100011011100000000110101110000111101110110000011011000" when "0001000000",
   "00001111101110000001110110100100101111111110001010010001010011110010001011" when "0001000001",
   "00001111111111000011010010000100110101011100100110000000010001100100110000" when "0001000010",
   "00001111111111000011010010000100110101011100100110000000010001100100110000" when "0001000011",
   "00010000010000000101110110000101111001110100010001000100011100000001011101" when "0001000100",
   "00010000100001001001100010110001100111100011101000000110100010001010010000" when "0001000101",
   "00010000110010001110011000010001101011000100111000010110110101000000010011" when "0001000110",
   "00010001000011010100010110101111110010101110100000110000100101101101011111" when "0001000111",
   "00010001010100011011011110010101101110110011110011001000100110101101111100" when "0001001000",
   "00010001100101100011101111001101010001100101010101100110110100010101010100" when "0001001001",
   "00010001110110101101001001100000001111010001100100001011001001001101100110" when "0001001010",
   "00010001110110101101001001100000001111010001100100001011001001001101100110" when "0001001011",
   "00010010000111110111101101011000011110000101010010011101100011001111110000" when "0001001100",
   "00010010011001000011011010111111110110001100001101101001011101011000000101" when "0001001101",
   "00010010101010010000010010100000010001110001011110100100100010111010100011" when "0001001110",
   "00010010111011011110010100000011101101000000001100000001000000111101101111" when "0001001111",
   "00010011001100101101011111110100000110000011111101001011011010100100101011" when "0001010000",
   "00010011011101111101110101111011011101001001011100010100000100010010100100" when "0001010001",
   "00010011011101111101110101111011011101001001011100010100000100010010100100" when "0001010010",
   "00010011101111001111010110100011110100011110111001100100001011110101001100" when "0001010011",
   "00010100000000100010000001110111010000010100101101111110110000100101010101" when "0001010100",
   "00010100010001110101110111111111110110111101111110101101010001101110100011" when "0001010101",
   "00010100100011001010111001000111110000110001000000011000010110110010000010" when "0001010110",
   "00010100110100100001000101011001001000000111111010101100010111011010011111" when "0001010111",
   "00010101000101111000011100111110001001100001001100001010000111011001011001" when "0001011000",
   "00010101000101111000011100111110001001100001001100001010000111011001011001" when "0001011001",
   "00010101010111010001000000000001000011100000001110000011101011101000000110" when "0001011010",
   "00010101101000101010101110101100000110101101111000100101011101001001111010" when "0001011011",
   "00010101111010000101101001001001100101111001000111001011011111001110000111" when "0001011100",
   "00010110001011100001101111100011110101110111011101000011001101010100000010" when "0001011101",
   "00010110011100111111000010000101001101100101101001111001100110010100110010" when "0001011110",
   "00010110011100111111000010000101001101100101101001111001100110010100110010" when "0001011111",
   "00010110101110011101100000111000000110001000001110110101111001111001100000" when "0001100000",
   "00010110111111111101001100000110111010101100000011100000111101000110110101" when "0001100001",
   "00010111010001011110000011111100001000100110111011011001001011101001001000" when "0001100010",
   "00010111100011000000001000100010001111011000001011010011011010101111001010" when "0001100011",
   "00010111110100100011011010000011110000101001001111001000100011000011111010" when "0001100100",
   "00010111110100100011011010000011110000101001001111001000100011000011111010" when "0001100101",
   "00011000000110000111111000101011010000001110001111110000000110111001111101" when "0001100110",
   "00011000010111101101100100100011010100000110101001000111111001111110011010" when "0001100111",
   "00011000101001010100011101110110100100011101110000101000110000001010111110" when "0001101000",
   "00011000111010111100100100101111101011101011011011101000011000110010000011" when "0001101001",
   "00011001001100100101111001011001010110010100100110001000101011100001110110" when "0001101010",
   "00011001001100100101111001011001010110010100100110001000101011100001110110" when "0001101011",
   "00011001011110010000011011111110010011001011111001110100001100111110100011" when "0001101100",
   "00011001101111111100001100101001010011010010010101001000001111110110000110" when "0001101101",
   "00011010000001101001001011100101001001110111110010101100011000110010011011" when "0001101110",
   "00011010010011010111011000111100101100011011110000110111101010010010100011" when "0001101111",
   "00011010010011010111011000111100101100011011110000110111101010010010100011" when "0001110000",
   "00011010100101000110110100111010110010101101111001100011011110010100110000" when "0001110001",
   "00011010110110110111011111101010010110101110101010001100010011011111011001" when "0001110010",
   "00011011001000101001011001010110010100101111111100000000010011011000100011" when "0001110011",
   "00011011011010011100100010001001101011010101101100011011110111111111010100" when "0001110100",
   "00011011101100010000111010001111011011010110100101110100010101111100101011" when "0001110101",
   "00011011101100010000111010001111011011010110100101110100010101111100101011" when "0001110110",
   "00011011111110000110100001110010100111111100101000010000110001100100011011" when "0001110111",
   "00011100001111111101011000111110010110100101110010110001000100100001110100" when "0001111000",
   "00011100100001110101011111111101101111000100101100100011011010001110001101" when "0001111001",
   "00011100110011101110110110111011111011100001001110101000001000110011000000" when "0001111010",
   "00011100110011101110110110111011111011100001001110101000001000110011000000" when "0001111011",
   "00011101000101101001011110000100001000011001001101100100001100111011011000" when "0001111100",
   "00011101010111100101010101100001100100100001000011100010001110011100110000" when "0001111101",
   "00011101101001100010011101011111100001000100011010100010010100000000100000" when "0001111110",
   "00011101101001100010011101011111100001000100011010100010010100000000100000" when "0001111111",
   "00011101111011100000110110001001010001100110110110111000101011111011111011" when "0010000000",
   "00011110001101100000011111101010001100000100100001111011010000100111001101" when "0010000001",
   "00011110011111100001011010001101101000110010110100111110001110100110010001" when "0010000010",
   "00011110110001100011100101111111000010100001000100011111110010111010100000" when "0010000011",
   "00011110110001100011100101111111000010100001000100011111110010111010100000" when "0010000100",
   "00011111000011100111000011001001110110011001001011100011000111110110110001" when "0010000101",
   "00011111010101101011110001111001100100000000010111011010100110110010011111" when "0010000110",
   "00011111100111110001110010011001101101010111110011100001100101011100000011" when "0010000111",
   "00011111111001111001000100110101110110111101010101100101100101001101100001" when "0010001000",
   "00011111111001111001000100110101110110111101010101100101100101001101100001" when "0010001001",
   "00100000001100000001101001011001100111101100001001111111001011001010001110" when "0010001010",
   "00100000011110001011100000010000101000111101100000011010100111001111000110" when "0010001011",
   "00100000110000010110101001100110100110101001011000110000010001100010100001" when "0010001100",
   "00100000110000010110101001100110100110101001011000110000010001100010100001" when "0010001101",
   "00100001000010100011000101100111001111000111010000001101000100010100100000" when "0010001110",
   "00100001010100110000110100011110010011001110101110101010111001100010100100" when "0010001111",
   "00100001100110111111110110010111100110011000010100011001010010110110101100" when "0010010000",
   "00100001111001010000001011011110111110011110000111110110010010111011111001" when "0010010001",
   "00100001111001010000001011011110111110011110000111110110010010111011111001" when "0010010010",
   "00100010001011100001110100000000010011111100100011110111101111000110011100" when "0010010011",
   "00100010011101110100110000000111100001110011000110000101000000010001001110" when "0010010100",
   "00100010110000001001000000000000100101100100111101100001011010010101010010" when "0010010101",
   "00100010110000001001000000000000100101100100111101100001011010010101010010" when "0010010110",
   "00100011000010011110100011110111011111011001111001100111010001000100010111" when "0010010111",
   "00100011010100110101011011111000010001111110111001010011110001110010001000" when "0010011000",
   "00100011100111001101101000001111000010100110111010100011111000111100011100" when "0010011001",
   "00100011100111001101101000001111000010100110111010100011111000111100011100" when "0010011010",
   "00100011111001100111001001000111111001001011101010000010001011000101100101" when "0010011011",
   "00100100001100000001111110101111000000001110010011000101111000011000000011" when "0010011100",
   "00100100011110011110001001010000100100111000010000000011010010001110010000" when "0010011101",
   "00100100011110011110001001010000100100111000010000000011010010001110010000" when "0010011110",
   "00100100110000111011101000111000110110111011111010101101011010011101000100" when "0010011111",
   "00100101000011011010011101110100001000110101011101001001010011100011010110" when "0010100000",
   "00100101010101111010101000001110101111101011100010110010111001100100101111" when "0010100001",
   "00100101010101111010101000001110101111101011100010110010111001100100101111" when "0010100010",
   "00100101101000011100001000010101000011010000001001110011101011011001100110" when "0010100011",
   "00100101111010111110111110010011011110000001010100101011001100000010000110" when "0010100100",
   "00100110001101100011001010010110011101001001111100001001100011101110001110" when "0010100101",
   "00100110001101100011001010010110011101001001111100001001100011101110001110" when "0010100110",
   "00100110100000001000101100101010100000100010100001011100001000110000100000" when "0010100111",
   "00100110110010101111100101011100001010110010000000101100010111110101000001" when "0010101000",
   "00100111000101010111110100111000000001001110100011110001000011111010101110" when "0010101001",
   "00100111000101010111110100111000000001001110100011110001000011111010101110" when "0010101010",
   "00100111011000000001011011001010101011111110010101010010000101110000110110" when "0010101011",
   "00100111101010101100011000100000110101111000010011111110110010111110000101" when "0010101100",
   "00100111101010101100011000100000110101111000010011111110110010111110000101" when "0010101101",
   "00100111111101011000101101000111001100100101000110010111000100111100000011" when "0010101110",
   "00101000010000000110011001001010100000011111101110100111010111110100111000" when "0010101111",
   "00101000100010110101011100110111100100110110011110110111101001110101100100" when "0010110000",
   "00101000100010110101011100110111100100110110011110110111101001110101100100" when "0010110001",
   "00101000110101100101111000011011001111101011101101101101100011001011111000" when "0010110010",
   "00101001001000010111101100000010011001110110101011000001101111001010101010" when "0010110011",
   "00101001011011001010110111111001111111000100010101001000101110110011110110" when "0010110100",
   "00101001011011001010110111111001111111000100010101001000101110110011110110" when "0010110101",
   "00101001101101111111011100001110111101111000001110001111001101101100000110" when "0010110110",
   "00101010000000110101011001001110010111101101010010001010000001011111111101" when "0010110111",
   "00101010000000110101011001001110010111101101010010001010000001011111111101" when "0010111000",
   "00101010010011101100101111000101010000110110101100011001111101000111001011" when "0010111001",
   "00101010100110100101011110000000110000100000101110100011011111110111001100" when "0010111010",
   "00101010111001011111100110001110000000110001100110111010101001111010011011" when "0010111011",
   "00101010111001011111100110001110000000110001100110111010101001111010011011" when "0010111100",
   "00101011001100011011000111111010001110101010010111100010111110100110100010" when "0010111101",
   "00101011011111011000000011010010101010000111101101100011111101110000010100" when "0010111110",
   "00101011011111011000000011010010101010000111101101100011111101110000010100" when "0010111111",
   "00101011110010010110011000100100100110000010111000110001111101000000110001" when "0011000000",
   "00101100000101010110000111111101011000010010100011101011101010010011011010" when "0011000001",
   "00101100011000010111010001101010011001101011101011101100100000101010110001" when "0011000010",
   "00101100011000010111010001101010011001101011101011101100100000101010110001" when "0011000011",
   "00101100101011011001110101111001000110000010011001110011111000101100101100" when "0011000100",
   "00101100111110011101110100110110111100001010111011100001011101111100111110" when "0011000101",
   "00101100111110011101110100110110111100001010111011100001011101111100111110" when "0011000110",
   "00101101010001100011001110110001011101111010011100000110110010110001100110" when "0011000111",
   "00101101100100101010000011110110010000000111111110001110001100000001010000" when "0011001000",
   "00101101110111110010010100010010111010101101010101110111001110010000110101" when "0011001001",
   "00101101110111110010010100010010111010101101010101110111001110010000110101" when "0011001010",
   "00101110001010111100000000010101001000101000000010101000110110001010110000" when "0011001011",
   "00101110011110000111001000001010100111111010001010011001010101101111001100" when "0011001100",
   "00101110011110000111001000001010100111111010001010011001010101101111001100" when "0011001101",
   "00101110110001010011101100000001001001101011010100001100010000010001110000" when "0011001110",
   "00101111000100100001101100000110100010001001100011100110011110111110010000" when "0011001111",
   "00101111000100100001101100000110100010001001100011100110011110111110010000" when "0011010000",
   "00101111010111110001001000101000101000101010010100011000101000000011010100" when "0011010001",
   "00101111101011000010000001110101010111101011010110011111110010100111010000" when "0011010010",
   "00101111101011000010000001110101010111101011010110011111110010100111010000" when "0011010011",
   "00101111111110010100010111111010101100110011101010011101000001010000001100" when "0011010100",
   "00110000010001101000001011000110101000110100011110000011011101101110011010" when "0011010101",
   "00110000100100111101011011100111001111101010001001011101011111111101010100" when "0011010110",
   "00110000100100111101011011100111001111101010001001011101011111111101010100" when "0011010111",
   "00110000111000010100001001101010101000011101001100101000111010110100001100" when "0011011000",
   "00110001001011101100010101011110111101100011001101001010011001000110010000" when "0011011001",
   "00110001001011101100010101011110111101100011001101001010011001000110010000" when "0011011010",
   "00110001011111000101111111010010011100011111110100011000010101010110101010" when "0011011011",
   "00110001110010100001000111010011010110000101101101111101010111001010101101" when "0011011100",
   "00110001110010100001000111010011010110000101101101111101010111001010101101" when "0011011101",
   "00110010000101111101101101101111111110010111100110110010100000101010001001" when "0011011110",
   "00110010011001011011110010110110101100101001001100010001010111000011101011" when "0011011111",
   "00110010011001011011110010110110101100101001001100010001010111000011101011" when "0011100000",
   "00110010101100111011010110110101111011100000001011111110010001010000101100" when "0011100001",
   "00110011000000011100011001111100001000110101010011101010110111011001111010" when "0011100010",
   "00110011000000011100011001111100001000110101010011101010110111011001111010" when "0011100011",
   "00110011010011111110111100010111110101110101010001110000111110100011111100" when "0011100100",
   "00110011100111100010111110010111100111000001110110000110001011110001000011" when "0011100101",
   "00110011100111100010111110010111100111000001110110000110001011110001000011" when "0011100110",
   "00110011111011001000100000001010000100010010110011001000001001101011010001" when "0011100111",
   "00110100001110101111100001111101111000110110111111100001111100001111111111" when "0011101000",
   "00110100001110101111100001111101111000110110111111100001111100001111111111" when "0011101001",
   "00110100100010011000000100000001110011010101011000001010011101111100100000" when "0011101010",
   "00110100110110000010000110100100100101101110000010011100010010000000111111" when "0011101011",
   "00110100110110000010000110100100100101101110000010011100010010000000111111" when "0011101100",
   "00110101001001101101101001110101000101011011001111000110110111100101011111" when "0011101101",
   "00110101011101011010101110000010001011010010011101011001101001010011010100" when "0011101110",
   "00110101011101011010101110000010001011010010011101011001101001010011010100" when "0011101111",
   "00110101110001001001010011011010110011100101011110101000110101011010111001" when "0011110000",
   "00110110000100111001011010001101111110000011011010001100011010010101001000" when "0011110001",
   "00110110000100111001011010001101111110000011011010001100011010010101001000" when "0011110010",
   "00110110011000101011000010101010101101111001110001111001010011100101011001" when "0011110011",
   "00110110101100011110001101000000001001110101100110110101000011101000001111" when "0011110100",
   "00110110101100011110001101000000001001110101100110110101000011101000001111" when "0011110101",
   "00110111000000010010111001011101011100000100011110100100000110100000111100" when "0011110110",
   "00110111000000010010111001011101011100000100011110100100000110100000111100" when "0011110111",
   "00110111010100001001001000010001110010010101101000110010111001111111010001" when "0011111000",
   "00110111101000000000111001101100011101111011000101011010000111011101001101" when "0011111001",
   "00110111101000000000111001101100011101111011000101011010000111011101001101" when "0011111010",
   "00110111111011111010001101111100110011101010101010111101111100011011010000" when "0011111011",
   "00111000001111110101000101010010001011111111001101101000111110001000110101" when "0011111100",
   "00111000001111110101000101010010001011111111001101101000111110001000110101" when "0011111101",
   "00111000100011110001011111111100000010111001100110100010100101001101011000" when "0011111110",
   "00111000110111101111011110001001111000000001111011100001001110001101001110" when "0011111111",
   "00111000110111101111011110001001111000000001111011100001001110001101001110" when "0100000000",
   "00111001001011101111000000001011001110101000100111011000101100001101010010" when "0100000001",
   "00111001011111110000000110001111101101100111100010100100101010011110100011" when "0100000010",
   "00111001011111110000000110001111101101100111100010100100101010011110100011" when "0100000011",
   "00111001110011110010110000100110111111100011001100001111101010100010111100" when "0100000100",
   "00111001110011110010110000100110111111100011001100001111101010100010111100" when "0100000101",
   "00111010000111110110111111100000110010101011110011110110101100000011000101" when "0100000110",
   "00111010011011111100110011001100111000111110100011001001101011110100110010" when "0100000111",
   "00111010011011111100110011001100111000111110100011001001101011110100110010" when "0100001000",
   "00111010110000000100001011111011001000000110101000101001000111111001000001" when "0100001001",
   "00111011000100001101001001111011011001011110100010100000110101111111110111" when "0100001010",
   "00111011000100001101001001111011011001011110100010100000110101111111110111" when "0100001011",
   "00111011011000010111101101011101101010010001001010000000011010101000010010" when "0100001100",
   "00111011101100100011110110110001111011011010111111010001001110011001011001" when "0100001101",
   "00111011101100100011110110110001111011011010111111010001001110011001011001" when "0100001110",
   "00111100000000110001100110001000010001101011010101101010011111111010100100" when "0100001111",
   "00111100000000110001100110001000010001101011010101101010011111111010100100" when "0100010000",
   "00111100010101000000111011110000110101100101100000100011100000010111011110" when "0100010001",
   "00111100101001010001110111111011110011100010000000100100001001000100111011" when "0100010010",
   "00111100101001010001110111111011110011100010000000100100001001000100111011" when "0100010011",
   "00111100111101100100011010111001011011101111110001010100001000100011101110" when "0100010100",
   "00111101010001111000100100111010000010010101010111101001000101100110001110" when "0100010101",
   "00111101010001111000100100111010000010010101010111101001000101100110001110" when "0100010110",
   "00111101100110001110010110001101111111010010010000010011100111000101110000" when "0100010111",
   "00111101100110001110010110001101111111010010010000010011100111000101110000" when "0100011000",
   "00111101111010100101101111000101101110011111111111001011101111011101010101" when "0100011001",
   "00111110001110111110101111110001101111110011011110111100111010100110110100" when "0100011010",
   "00111110001110111110101111110001101111110011011110111100111010100110110100" when "0100011011",
   "00111110100011011001011000100010100110111110010001010001101101100000111000" when "0100011100",
   "00111110100011011001011000100010100110111110010001010001101101100000111000" when "0100011101",
   "00111110110111110101101001101000111011101111101111011111100110101011101010" when "0100011110",
   "00111111001100010011100011010101011001110110011011110010111110110011001010" when "0100011111",
   "00111111001100010011100011010101011001110110011011110010111110110011001010" when "0100100000",
   "00111111100000110011000101111000110001000001010010111011101001000110111100" when "0100100001",
   "00111111100000110011000101111000110001000001010010111011101001000110111100" when "0100100010",
   "00111111110101010100010001100011110101000000111110011010000011000110111100" when "0100100011",
   "01000000001001110111000110100111011101101001000111001101100011010110100010" when "0100100100",
   "01000000001001110111000110100111011101101001000111001101100011010110100010" when "0100100101",
   "01000000011110011011100101010100100110110001101001000011110111001111101100" when "0100100110",
   "01000000110011000001101101111100010000011000000110001001111111111000101010" when "0100100111",
   "01000000110011000001101101111100010000011000000110001001111111111000101010" when "0100101000",
   "01000001000111101001100000101111011110100000111011011110111110001000011010" when "0100101001",
   "01000001000111101001100000101111011110100000111011011110111110001000011010" when "0100101010",
   "01000001011100010010111101111111011001011000110101101000011110001110001111" when "0100101011",
   "01000001110000111110000101111101001101010110000110001001110011011011000110" when "0100101100",
   "01000001110000111110000101111101001101010110000110001001110011011011000110" when "0100101101",
   "01000010000101101010111000111010001010111001111001011101010100010011111101" when "0100101110",
   "01000010000101101010111000111010001010111001111001011101010100010011111101" when "0100101111",
   "01000010011010011001010111000111100110110001101101010000101000011110000110" when "0100110000",
   "01000010101111001001100000110110111001111000100111100011111000011111101010" when "0100110001",
   "01000010101111001001100000110110111001111000100111100011111000011111101010" when "0100110010",
   "01000011000011111011010110011001100001011000101110001100010001011000101100" when "0100110011",
   "01000011000011111011010110011001100001011000101110001100010001011000101100" when "0100110100",
   "01000011011000101110111000000000111110101100011110111010001100100010001000" when "0100110101",
   "01000011011000101110111000000000111110101100011110111010001100100010001000" when "0100110110",
   "01000011101101100100000101111110110111100000001000000011001101101010010111" when "0100110111",
   "01000100000010011011000000100100110101110011000001110000001000010001000000" when "0100111000",
   "01000100000010011011000000100100110101110011000001110000001000010001000000" when "0100111001",
   "01000100010111010011101000000100100111111001000111101111011110001100111000" when "0100111010",
   "01000100010111010011101000000100100111111001000111101111011110001100111000" when "0100111011",
   "01000100101100001101111100110000000000011100010011101100101001010010001010" when "0100111100",
   "01000101000001001001111110111000110110011101111000001100000001111000001001" when "0100111101",
   "01000101000001001001111110111000110110011101111000001100000001111000001001" when "0100111110",
   "01000101010110000111101110110001000101010111111100001100010100101001000000" when "0100111111",
   "01000101010110000111101110110001000101010111111100001100010100101001000000" when "0101000000",
   "01000101101011000111001100101010101100111110110111001101011001101111110000" when "0101000001",
   "01000101101011000111001100101010101100111110110111001101011001101111110000" when "0101000010",
   "01000110000000001000011000110111110001100010101101111101000000000011011110" when "0101000011",
   "01000110010101001011010011101010011011110000101111101001011110111001110110" when "0101000100",
   "01000110010101001011010011101010011011110000101111101001011110111001110110" when "0101000101",
   "01000110101010001111111101010100111000110100110011111011000001010100101100" when "0101000110",
   "01000110101010001111111101010100111000110100110011111011000001010100101100" when "0101000111",
   "01000110111111010110010110001001011010011010111001010011011101101010100010" when "0101001000",
   "01000110111111010110010110001001011010011010111001010011011101101010100010" when "0101001001",
   "01000111010100011110011110011010010110110000100100010101001100110011111000" when "0101001010",
   "01000111101001101000010110011010001000100110011111010001010100010010110001" when "0101001011",
   "01000111101001101000010110011010001000100110011111010001010100010010110001" when "0101001100",
   "01000111111110110011111110011011001111010001111010011101010110110101000101" when "0101001101",
   "01000111111110110011111110011011001111010001111010011101010110110101000101" when "0101001110",
   "01001000010100000001010110110000001110101110001101010000111110111101011101" when "0101001111",
   "01001000010100000001010110110000001110101110001101010000111110111101011101" when "0101010000",
   "01001000101001010000011111101011101111011110010111101011110111101001111110" when "0101010001",
   "01001000111110100001011001100000011110101110100100100100000110111011011110" when "0101010010",
   "01001000111110100001011001100000011110101110100100100100000110111011011110" when "0101010011",
   "01001001010011110100000100100001001110010101101100011101011110101100000100" when "0101010100",
   "01001001010011110100000100100001001110010101101100011101011110101100000100" when "0101010101",
   "01001001101001001000100001000000110100110110111001001001111000001110111110" when "0101010110",
   "01001001101001001000100001000000110100110110111001001001111000001110111110" when "0101010111",
   "01001001111110011110101111010010001101100011001001110011001110111111111110" when "0101011000",
   "01001010010011110110101111101000011000011010110111101111001111010100100011" when "0101011001",
   "01001010010011110110101111101000011000011010110111101111001111010100100011" when "0101011010",
   "01001010101001010000100010010110011010001111011011111101001110001101010101" when "0101011011",
   "01001010101001010000100010010110011010001111011011111101001110001101010101" when "0101011100",
   "01001010111110101100000111101111011100100100110101001110011111010010010100" when "0101011101",
   "01001010111110101100000111101111011100100100110101001110011111010010010100" when "0101011110",
   "01001011010100001001100000000110101101110011001110111001011110010001000110" when "0101011111",
   "01001011010100001001100000000110101101110011001110111001011110010001000110" when "0101100000",
   "01001011101001101000101011101111100001001000101000011000000001100000100101" when "0101100001",
   "01001011111111001001101010111101001110101010011101010001001011011010110000" when "0101100010",
   "01001011111111001001101010111101001110101010011101010001001011011010110000" when "0101100011",
   "01001100010100101100011110000011010011010111001110001110110000101001011010" when "0101100100",
   "01001100010100101100011110000011010011010111001110001110110000101001011010" when "0101100101",
   "01001100101010010001000101010101010001001000001010011111001001010000001010" when "0101100110",
   "01001100101010010001000101010101010001001000001010011111001001010000001010" when "0101100111",
   "01001100111111110111100001000110101110110010111010000011100011001010101010" when "0101101000",
   "01001100111111110111100001000110101110110010111010000011100011001010101010" when "0101101001",
   "01001101010101011111110001101011011000001011001000101011001100100011101101" when "0101101010",
   "01001101010101011111110001101011011000001011001000101011001100100011101101" when "0101101011",
   "01001101101011001001110111010110111110000100010001011011101100110110110001" when "0101101100",
   "01001110000000110101110010011101010110010011001011000111000011011011011000" when "0101101101",
   "01001110000000110101110010011101010110010011001011000111000011011011011000" when "0101101110",
   "01001110010110100011100011010010011011101111110101001111100011000111010101" when "0101101111",
   "01001110010110100011100011010010011011101111110101001111100011000111010101" when "0101110000",
   "01001110101100010011001010001010001110010111000101111010000010000010001000" when "0101110001",
   "01001110101100010011001010001010001110010111000101111010000010000010001000" when "0101110010",
   "01001111000010000100100111011000110011001100011000001110110101010010110110" when "0101110011",
   "01001111000010000100100111011000110011001100011000001110110101010010110110" when "0101110100",
   "01001111010111110111111011010010010100011011011011101001110000011110101011" when "0101110101",
   "01001111010111110111111011010010010100011011011011101001110000011110101011" when "0101110110",
   "01001111101101101101000110001011000001011010000011111001100000111101011010" when "0101110111",
   "01010000000011100100001000010111001110101001111001101110111101010111010001" when "0101111000",
   "01010000000011100100001000010111001110101001111001101110111101010111010001" when "0101111001",
   "01010000011001011101000010001011010101111010001100011100100001101101110110" when "0101111010",
   "01010000011001011101000010001011010101111010001100011100100001101101110110" when "0101111011",
   "01010000101111010111110011111011110110001001100100000110010001000000111110" when "0101111100",
   "01010000101111010111110011111011110110001001100100000110010001000000111110" when "0101111101",
   "01010001000101010100011101111101010011100111110100100010110101001110110110" when "0101111110",
   "01010001000101010100011101111101010011100111110100100010110101001110110110" when "0101111111",
   "01010001011011010011000000100100010111110111110001001101110110111110001100" when "0110000000",
   "01010001011011010011000000100100010111110111110001001101110110111110001100" when "0110000001",
   "01010001110001010011011100000101110001110001000001101100000110001111101101" when "0110000010",
   "01010001110001010011011100000101110001110001000001101100000110001111101101" when "0110000011",
   "01010010000111010101110000110110010101100001110111000001101110000100011010" when "0110000100",
   "01010010000111010101110000110110010101100001110111000001101110000100011010" when "0110000101",
   "01010010011101011001111111001010111100110001000001111011001100110100110110" when "0110000110",
   "01010010011101011001111111001010111100110001000001111011001100110100110110" when "0110000111",
   "01010010110011100000000111011000100110011111101001101001001011100101111111" when "0110001000",
   "01010011001001101000001001110100010111001011000011101111101110110111001010" when "0110001001",
   "01010011001001101000001001110100010111001011000011101111101110110111001010" when "0110001010",
   "01010011011111110010000110110011011000101110101100101001011011010101111000" when "0110001011",
   "01010011011111110010000110110011011000101110101100101001011011010101111000" when "0110001100",
   "01010011110101111101111110101010111010100110000000111110101001110011010011" when "0110001101",
   "01010011110101111101111110101010111010100110000000111110101001110011010011" when "0110001110",
   "01010100001100001011110001110000010001101110010111110001100101001000000110" when "0110001111",
   "01010100001100001011110001110000010001101110010111110001100101001000000110" when "0110010000",
   "01010100100010011011100000011000111000101000111101011111001110000100000011" when "0110010001",
   "01010100100010011011100000011000111000101000111101011111001110000100000011" when "0110010010",
   "01010100111000101101001010111010001111011100101111110110000000010111001000" when "0110010011",
   "01010100111000101101001010111010001111011100101111110110000000010111001000" when "0110010100",
   "01010101001111000000110001101001111011111000011010100010010101010011000000" when "0110010101",
   "01010101001111000000110001101001111011111000011010100010010101010011000000" when "0110010110",
   "01010101100101010110010100111101101001010100010100110001011111110100101100" when "0110010111",
   "01010101100101010110010100111101101001010100010100110001011111110100101100" when "0110011000",
   "01010101111011101101110101001011001000110100011111101011011110110111101110" when "0110011001",
   "01010101111011101101110101001011001000110100011111101011011110110111101110" when "0110011010",
   "01010110010010000111010010101000010001001010100101100100000010100101100010" when "0110011011",
   "01010110010010000111010010101000010001001010100101100100000010100101100010" when "0110011100",
   "01010110101000100010101101101010111110110111111010000011100001100100111110" when "0110011101",
   "01010110101000100010101101101010111110110111111010000011100001100100111110" when "0110011110",
   "01010110111111000000000110101001010100001111011011000111111011100000101001" when "0110011111",
   "01010110111111000000000110101001010100001111011011000111111011100000101001" when "0110100000",
   "01010111010101011111011101111001011001010111110010111110100110101011111100" when "0110100001",
   "01010111010101011111011101111001011001010111110010111110100110101011111100" when "0110100010",
   "01010111101100000000110011110001011100001101011010110111000110100001001000" when "0110100011",
   "01010111101100000000110011110001011100001101011010110111000110100001001000" when "0110100100",
   "01011000000010100100001000100111110000100100011110101111101001000101110111" when "0110100101",
   "01011000000010100100001000100111110000100100011110101111101001000101110111" when "0110100110",
   "01011000011001001001011100110010110000001011000001111011101010010101000000" when "0110100111",
   "01011000011001001001011100110010110000001011000001111011101010010101000000" when "0110101000",
   "01011000101111110000110000101000111010101011000100100100111011100000110010" when "0110101001",
   "01011000101111110000110000101000111010101011000100100100111011100000110010" when "0110101010",
   "01011001000110011010000100100000110101101100101010000111101110010010010111" when "0110101011",
   "01011001000110011010000100100000110101101100101010000111101110010010010111" when "0110101100",
   "01011001011101000101011000110001001100111000000000101010100010011111101010" when "0110101101",
   "01011001011101000101011000110001001100111000000000101010100010011111101010" when "0110101110",
   "01011001110011110010101101110000110001110111101001010001110110100011101010" when "0110101111",
   "01011001110011110010101101110000110001110111101001010001110110100011101010" when "0110110000",
   "01011010001010100010000011110110011100011010100001010000011010011001001110" when "0110110001",
   "01011010001010100010000011110110011100011010100001010000011010011001001110" when "0110110010",
   "01011010100001010011011011011001001010010110001100010100100101001100001010" when "0110110011",
   "01011010100001010011011011011001001010010110001100010100100101001100001010" when "0110110100",
   "01011010111000000110110100101111111111101000111111110011001110101000011010" when "0110110101",
   "01011010111000000110110100101111111111101000111111110011001110101000011010" when "0110110110",
   "01011011001110111100010000010010000110011100001110110000101100100100010010" when "0110110111",
   "01011011001110111100010000010010000110011100001110110000101100100100010010" when "0110111000",
   "01011011100101110011101110010110101111000110010111001000010110010101111100" when "0110111001",
   "01011011100101110011101110010110101111000110010111001000010110010101111100" when "0110111010",
   "01011011111100101101001111010101010000001101001111110011001111011010100000" when "0110111011",
   "01011011111100101101001111010101010000001101001111110011001111011010100000" when "0110111100",
   "01011100010011101000110011100101000110101000010111101110011011001001100010" when "0110111101",
   "01011100010011101000110011100101000110101000010111101110011011001001100010" when "0110111110",
   "01011100101010100110011011011101110101100011000110000001011100000100110010" when "0110111111",
   "01011100101010100110011011011101110101100011000110000001011100000100110010" when "0111000000",
   "01011101000001100110000111010111000110011110111011000101100001001010010100" when "0111000001",
   "01011101000001100110000111010111000110011110111011000101100001001010010100" when "0111000010",
   "01011101011000100111110111101000101001010101110010101110000100000100001010" when "0111000011",
   "01011101011000100111110111101000101001010101110010101110000100000100001010" when "0111000100",
   "01011101101111101011101100101010010100011100010111010010111011100111001010" when "0111000101",
   "01011101101111101011101100101010010100011100010111010010111011100111001010" when "0111000110",
   "01011110000110110001100110110100000100100100010101111101000110001000101000" when "0111000111",
   "01011110000110110001100110110100000100100100010101111101000110001000101000" when "0111001000",
   "01011110000110110001100110110100000100100100010101111101000110001000101000" when "0111001001",
   "01011110011101111001100110011101111100111110110011110110001111101001011110" when "0111001010",
   "01011110011101111001100110011101111100111110110011110110001111101001011110" when "0111001011",
   "01011110110101000011101100000000000111011110100100011011111000001011011000" when "0111001100",
   "01011110110101000011101100000000000111011110100100011011111000001011011000" when "0111001101",
   "01011111001100001111110111110010110100011010100000110110011110111100100000" when "0111001110",
   "01011111001100001111110111110010110100011010100000110110011110111100100000" when "0111001111",
   "01011111100011011110001010001110011010110000000000010101010111011101000110" when "0111010000",
   "01011111100011011110001010001110011010110000000000010101010111011101000110" when "0111010001",
   "01011111111010101110100011101011011000000101010001101111101101111001110000" when "0111010010",
   "01011111111010101110100011101011011000000101010001101111101101111001110000" when "0111010011",
   "01100000010010000001000100100010010000101011110110001011100000101101011010" when "0111010100",
   "01100000010010000001000100100010010000101011110110001011100000101101011010" when "0111010101",
   "01100000101001010101101101001011101111100010111100101010110101010101110100" when "0111010110",
   "01100000101001010101101101001011101111100010111100101010110101010101110100" when "0111010111",
   "01100001000000101100011110000000100110011001111111000000001110111101110111" when "0111011000",
   "01100001000000101100011110000000100110011001111111000000001110111101110111" when "0111011001",
   "01100001011000000101010111011001101101110010111111101010101101111001100110" when "0111011010",
   "01100001011000000101010111011001101101110010111111101010101101111001100110" when "0111011011",
   "01100001011000000101010111011001101101110010111111101010101101111001100110" when "0111011100",
   "01100001101111100000011001110000000101000101001000111001111111001000111100" when "0111011101",
   "01100001101111100000011001110000000101000101001000111001111111001000111100" when "0111011110",
   "01100010000110111101100101011100110010011111001100111011100011101111000001" when "0111011111",
   "01100010000110111101100101011100110010011111001100111011100011101111000001" when "0111100000",
   "01100010011110011100111010111001000011001010000111010001011000000110000100" when "0111100001",
   "01100010011110011100111010111001000011001010000111010001011000000110000100" when "0111100010",
   "01100010110101111110011010011110001011001011011111010010100011110000110100" when "0111100011",
   "01100010110101111110011010011110001011001011011111010010100011110000110100" when "0111100100",
   "01100011001101100010000100100101100101101000001011110110111010100101011010" when "0111100101",
   "01100011001101100010000100100101100101101000001011110110111010100101011010" when "0111100110",
   "01100011100101000111111001101000110100100110111000001101111000100111011001" when "0111100111",
   "01100011100101000111111001101000110100100110111000001101111000100111011001" when "0111101000",
   "01100011100101000111111001101000110100100110111000001101111000100111011001" when "0111101001",
   "01100011111100101111111010000001100001010010101010000001100010100001100010" when "0111101010",
   "01100011111100101111111010000001100001010010101010000001100010100001100010" when "0111101011",
   "01100100010100011010000110001001011011111101101000100110010100101011010001" when "0111101100",
   "01100100010100011010000110001001011011111101101000100110010100101011010001" when "0111101101",
   "01100100101100000110011110011010011100000011100101011000001011100000011101" when "0111101110",
   "01100100101100000110011110011010011100000011100101011000001011100000011101" when "0111101111",
   "01100101000011110101000011001110100000001100100101100101110000001110010010" when "0111110000",
   "01100101000011110101000011001110100000001100100101100101110000001110010010" when "0111110001",
   "01100101011011100101110100111111101110001111101101001010010101010011111010" when "0111110010",
   "01100101011011100101110100111111101110001111101101001010010101010011111010" when "0111110011",
   "01100101011011100101110100111111101110001111101101001010010101010011111010" when "0111110100",
   "01100101110011011000110100001000010011010101101010110111001110110001011011" when "0111110101",
   "01100101110011011000110100001000010011010101101010110111001110110001011011" when "0111110110",
   "01100110001011001110000001000010100011111011100101101101010010011101001100" when "0111110111",
   "01100110001011001110000001000010100011111011100101101101010010011101001100" when "0111111000",
   "01100110100011000101011100001000111011110101101011100111001101010011010101" when "0111111001",
   "01100110100011000101011100001000111011110101101011100111001101010011010101" when "0111111010",
   "01100110111010111111000101110101111110010010000001010101011010110001110000" when "0111111011",
   "01100110111010111111000101110101111110010010000001010101011010110001110000" when "0111111100",
   "01100110111010111111000101110101111110010010000001010101011010110001110000" when "0111111101",
   "01100111010010111010111110100100010101111011010011101100001100001111011110" when "0111111110",
   "01100111010010111010111110100100010101111011010011101100001100001111011110" when "0111111111",
   "10110110001110010111100110110111000000011110101100001011000011100000101000" when "1000000000",
   "10110110011010010111100000110111001100011110011101001011011101111001100100" when "1000000001",
   "10110110100110010111111110111000100000100010011100011000010000111101110111" when "1000000010",
   "10110110110010011001000000111110010101000100000000011101110101111000000100" when "1000000011",
   "10110110111110011010100111001100000010111010111111110000000000001100111000" when "1000000100",
   "10110111001010011100110001100101000011011101110101111000111011010000011000" when "1000000101",
   "10110111001010011100110001100101000011011101110101111000111011010000011000" when "1000000110",
   "10110111010110011111100000001100110000100001101001101001011101101111011000" when "1000000111",
   "10110111100010100010110011000110100100011010010010101010110100000100110110" when "1000001000",
   "10110111101110100110101010010101111001111010011111010001100001110100011000" when "1000001001",
   "10110111111010101011000101111110001100010011111010010001111010100001111010" when "1000001010",
   "10111000000110110000000110000010110111010111010000110101110010011111111000" when "1000001011",
   "10111000010010110101101010100111010111010100011000010011100111101100001010" when "1000001100",
   "10111000011110111011110011101111001000111010010100000111000011010101011001" when "1000001101",
   "10111000011110111011110011101111001000111010010100000111000011010101011001" when "1000001110",
   "10111000101011000010100001011101101001010111011011101010110100100001011101" when "1000001111",
   "10111000110111001001110011110110010110011001100000010100000100001110010111" when "1000010000",
   "10111001000011010001101010111100101110001101110011001111000011000111010010" when "1000010001",
   "10111001001111011010000110110100001111100001001011011101010001100110110111" when "1000010010",
   "10111001011011100011000111100000011001100000001011110101000010100000110010" when "1000010011",
   "10111001100111101100101101000100101011110111001001000010011000101100001100" when "1000010100",
   "10111001110011110110110111100100100110110010001111101001100000001001000011" when "1000010101",
   "10111001110011110110110111100100100110110010001111101001100000001001000011" when "1000010110",
   "10111010000000000001100111000011101010111101101010001010100010111010011101" when "1000010111",
   "10111010001100001100111011100101011001100101100111000110111010010000000001" when "1000011000",
   "10111010011000011000110101001101010100010110011111000111111100011000110100" when "1000011001",
   "10111010100100100101010011111110111101011100111011000111000111011010010100" when "1000011010",
   "10111010110000110010010111111101110111100101111010010111101001100101111000" when "1000011011",
   "10111010111101000000000001001101100101111110111000110001100111100111101001" when "1000011100",
   "10111010111101000000000001001101100101111110111000110001100111100111101001" when "1000011101",
   "10111011001001001110001111110001101100010101110100111110100001001001101000" when "1000011110",
   "10111011010101011101000011101101101110111001010110100111010100000110000101" when "1000011111",
   "10111011100001101100011101000101010010011000110100100011111111000100100000" when "1000100000",
   "10111011101101111100011011111011111100000100011011001100100011011100001010" when "1000100001",
   "10111011111010001101000000010101010001101101010010101011100111011000000110" when "1000100010",
   "10111100000110011110001010010100111001100101100101010010011000010111111100" when "1000100011",
   "10111100000110011110001010010100111001100101100101010010011000010111111100" when "1000100100",
   "10111100010010101111111001111110011010100000100101101110001110101001010000" when "1000100101",
   "10111100011111000010001111010101011011110010110101011111110001110101100010" when "1000100110",
   "10111100101011010101001010011101100101010010001011010011011111100000100111" when "1000100111",
   "10111100110111101000101011011010011111010101111001011011110011110100000000" when "1000101000",
   "10111101000011111100110010001111110010110110110100001100110100110011001110" when "1000101001",
   "10111101010000010001011111000001001001001111011000011001100000110101101110" when "1000101010",
   "10111101010000010001011111000001001001001111011000011001100000110101101110" when "1000101011",
   "10111101011100100110110001110010001100011011110001110010100000100011000000" when "1000101100",
   "10111101101000111100101010100110100110111010000001100110011100101101111110" when "1000101101",
   "10111101110101010011001001100010000011101010000101000011111000101011111101" when "1000101110",
   "10111110000001101010001110101000001110001101111011111100110001100100111101" when "1000101111",
   "10111110001110000001111001111100110010101001101111001011100010111010010000" when "1000110000",
   "10111110001110000001111001111100110010101001101111001011100010111010010000" when "1000110001",
   "10111110011010011010001011100011011101100011110111011001110001000000100110" when "1000110010",
   "10111110100110110011000011011111111100000101000011101000011001101011110100" when "1000110011",
   "10111110110011001100100001110101111011111000011111111001101011101001010001" when "1000110100",
   "10111110111111100110100110101001001011001011111011111100100101000111011000" when "1000110101",
   "10111111001100000001010001111101011000101111110001111001111010000111110110" when "1000110110",
   "10111111001100000001010001111101011000101111110001111001111010000111110110" when "1000110111",
   "10111111011000011100100011110110010011110111001101000011000010111011000110" when "1000111000",
   "10111111100100111000011100010111101100011000010000100010010011000011001101" when "1000111001",
   "10111111110001010100111011100101010010101011111110001100111001011100101011" when "1000111010",
   "10111111111101110010000001100010110111101110011101010110101010001011111101" when "1000111011",
   "10111111111101110010000001100010110111101110011101010110101010001011111101" when "1000111100",
   "11000000001010001111101110010100001100111111000001100111010010001110011010" when "1000111101",
   "11000000010110101110000001111101000100100000010001110001010101101101110011" when "1000111110",
   "11000000100011001100111100100001010000111000001110101010111001010101010110" when "1000111111",
   "11000000101111101100011110000100100101010000011010000111110111000111111011" when "1001000000",
   "11000000111100001100100110101010110101010101111101110101111111010110101001" when "1001000001",
   "11000000111100001100100110101010110101010101111101110101111111010110101001" when "1001000010",
   "11000001001000101101010110010111110101011001110010011010100101110111101011" when "1001000011",
   "11000001010101001110101101001111011010010000100110010001111100011101000001" when "1001000100",
   "11000001100001110000101011010101011001010011000100110000011010101011011001" when "1001000101",
   "11000001101110010011010000101101101000011101111101000101010011110001010000" when "1001000110",
   "11000001101110010011010000101101101000011101111101000101010011110001010000" when "1001000111",
   "11000001111010110110011101011011111110010010001001011111011010111110011100" when "1001001000",
   "11000010000111011010010001100100010001110100110110010011010110111100111001" when "1001001001",
   "11000010010011111110101101001010011010101111101001000011100100101011001000" when "1001001010",
   "11000010100000100011110000010010010001010000100111101010001010011001100010" when "1001001011",
   "11000010101101001001011010111111101110001010011111100100011011001011001110" when "1001001100",
   "11000010101101001001011010111111101110001010011111100100011011001011001110" when "1001001101",
   "11000010111001101111101101010110101010110100101101000000001011011100000010" when "1001001110",
   "11000011000110010110100111011011000001001011100010001010110111001100110010" when "1001001111",
   "11000011010010111110001001010000101011110000001110100010011010010111101000" when "1001010000",
   "11000011011111100110010010111011100101101001000110000111111011101110000010" when "1001010001",
   "11000011011111100110010010111011100101101001000110000111111011101110000010" when "1001010010",
   "11000011101100001111000100011111101010100001101000110100001011000010101100" when "1001010011",
   "11000011111000111000011110000000110110101010101001101101110011000000111111" when "1001010100",
   "11000100000101100010011111100011000110111010010110100001011111010100111101" when "1001010101",
   "11000100010010001101001001001010011000101100011110111011110111100101110001" when "1001010110",
   "11000100010010001101001001001010011000101100011110111011110111100101110001" when "1001010111",
   "11000100011110111000011010111010101010000010011100000101001111100101100111" when "1001011000",
   "11000100101011100100010100110111111001100011010111111111001101011001111101" when "1001011001",
   "11000100111000010000110111000110000110011100010101000100000101111111000100" when "1001011010",
   "11000101000100111110000001101001010000100000010101101000010000101010001011" when "1001011011",
   "11000101000100111110000001101001010000100000010101101000010000101010001011" when "1001011100",
   "11000101010001101011110100100101011000001000100011011101010010001101111000" when "1001011101",
   "11000101011110011010001111111110011110010100010111010111000000000011111110" when "1001011110",
   "11000101101011001001010011111000100100101001100000110010011100000001001010" when "1001011111",
   "11000101101011001001010011111000100100101001100000110010011100000001001010" when "1001100000",
   "11000101110111111001000000010111101101010100001101011110101001010110010000" when "1001100001",
   "11000110000100101001010101011111111011000111010001000111011011100011001100" when "1001100010",
   "11000110010001011010010011010101010001011100001101000001111111100000011010" when "1001100011",
   "11000110011110001011111001111011110100010011010111111011011111100011001011" when "1001100100",
   "11000110011110001011111001111011110100010011010111111011011111100011001011" when "1001100101",
   "11000110101010111110001001010111101000010100000101101001100011000001100011" when "1001100110",
   "11000110110111110001000001101100110010101100101110111100101001111011010001" when "1001100111",
   "11000111000100100100100010111111011001010010111001010100100101001100100110" when "1001101000",
   "11000111010001011000101101010011100010100011011110110110101100010000100110" when "1001101001",
   "11000111010001011000101101010011100010100011011110110110101100010000100110" when "1001101010",
   "11000111011110001101100000101101010101100010110110000110010000011000101101" when "1001101011",
   "11000111101011000010111101010000111001111100111001111110101110011110111110" when "1001101100",
   "11000111110111111001000011000010011000000101010001101111111111111001101000" when "1001101101",
   "11000111110111111001000011000010011000000101010001101111111111111001101000" when "1001101110",
   "11001000000100101111110010000101111000110111011000111100101010110101110000" when "1001101111",
   "11001000010001100111001010011111100101110110100111011010010010111111110111" when "1001110000",
   "11001000011110011111001100010011101001001110011001010011101011000000110010" when "1001110001",
   "11001000011110011111001100010011101001001110011001010011101011000000110010" when "1001110010",
   "11001000101011010111110111100110001101110010010111001101000111010110000100" when "1001110011",
   "11001000111000010001001100011011011110111110011110001010110011001100111000" when "1001110100",
   "11001001000101001011001010110111101000110111000111111001001000000110100011" when "1001110101",
   "11001001010010000101110010111110111000001001010010110111001000101110110000" when "1001110110",
   "11001001010010000101110010111110111000001001010010110111001000101110110000" when "1001110111",
   "11001001011111000001000100110101011010001010101010100010111111101010100110" when "1001111000",
   "11001001101011111101000000011111011100111001101111101000100010101001000010" when "1001111001",
   "11001001111000111001100110000001001110111110000000010001111010111100011100" when "1001111010",
   "11001001111000111001100110000001001110111110000000010001111010111100011100" when "1001111011",
   "11001010000101110110110101011110111111101000000000011010010011100110001101" when "1001111100",
   "11001010010010110100101110111100111110110001100010000010101101111100100000" when "1001111101",
   "11001010011111110011010010011111011100111101101101101000111101010011100110" when "1001111110",
   "11001010011111110011010010011111011100111101101101101000111101010011100110" when "1001111111",
   "11001010101100110010100000001010101011011001001010100000101010010011011010" when "1010000000",
   "11001010111001110010011000000010111011111010000111001110011110100011000100" when "1010000001",
   "11001011000110110010111010001100100001000000100010000101011001010011011110" when "1010000010",
   "11001011000110110010111010001100100001000000100010000101011001010011011110" when "1010000011",
   "11001011010011110100000110101011101101110110010001100110001101110011011000" when "1010000100",
   "11001011100000110101111101100100110110001111001101000001001011110110010011" when "1010000101",
   "11001011101101111000011110111100001110101001010100111001110011011001001000" when "1010000110",
   "11001011101101111000011110111100001110101001010100111001110011011001001000" when "1010000111",
   "11001011111010111011101010110110001100001100111011101100110011101110011010" when "1010001000",
   "11001100000111111111100001010111000100101100101110011000010110111101101000" when "1010001001",
   "11001100010101000100000010100011001110100101111101000110011010011111110001" when "1010001010",
   "11001100010101000100000010100011001110100101111101000110011010011111110001" when "1010001011",
   "11001100100010001001001110011111000001000000100011111001010101000101000100" when "1010001100",
   "11001100101111001111000101001110110011101111010011011010101011001110111000" when "1010001101",
   "11001100111100010101100110110110111111001111111001101100010010101001101100" when "1010001110",
   "11001100111100010101100110110110111111001111111001101100010010101001101100" when "1010001111",
   "11001101001001011100110011011011111100101011001010111011100101010011000110" when "1010010000",
   "11001101010110100100101011000010000101110101001010010111000100110111110110" when "1010010001",
   "11001101100011101101001101101101110101001101010011000110001111010110101001" when "1010010010",
   "11001101100011101101001101101101110101001101010011000110001111010110101001" when "1010010011",
   "11001101110000110110011011100011100101111110100001000011100101010100001000" when "1010010100",
   "11001101111110000000010100100111110011111111011001111001000010101101010000" when "1010010101",
   "11001110001011001010111000111110111011110010010101111110101010110100111011" when "1010010110",
   "11001110001011001010111000111110111011110010010101111110101010110100111011" when "1010010111",
   "11001110011000010110001000101101011010100101101001011011101000001010101001" when "1010011000",
   "11001110100101100010000011110111101110010011101101001001100000110111110000" when "1010011001",
   "11001110110010101110101010100010010101100011000111111010000000100001001011" when "1010011010",
   "11001110110010101110101010100010010101100011000111111010000000100001001011" when "1010011011",
   "11001110111111111011111100110001101111100110110111011110110111111100000000" when "1010011100",
   "11001111001101001001111010101010011100011110011001110100010011110011010011" when "1010011101",
   "11001111011010011000100100010000111100110101110110001101101010101101111101" when "1010011110",
   "11001111011010011000100100010000111100110101110110001101101010101101111101" when "1010011111",
   "11001111100111100111111001101001110010000110000110100100100011100011100100" when "1010100000",
   "11001111110100110111111010111001011110010101000000101010010100101111100100" when "1010100001",
   "11001111110100110111111010111001011110010101000000101010010100101111100100" when "1010100010",
   "11010000000010001000101000000100100100010101011111011011111101010010010010" when "1010100011",
   "11010000001111011010000001001111100111100111101100011000011000001111100010" when "1010100100",
   "11010000011100101100000110011111001100011001001000111001001011011011001100" when "1010100101",
   "11010000011100101100000110011111001100011001001000111001001011011011001100" when "1010100110",
   "11010000101001111110110111110111110111100100110111101101110010000011100101" when "1010100111",
   "11010000110111010010010101011110001110110011100110011001000100001010110010" when "1010101000",
   "11010000110111010010010101011110001110110011100110011001000100001010110010" when "1010101001",
   "11010001000100100110011111010110111000011011110110110001011011011111100110" when "1010101010",
   "11010001010001111011010101100110011011100010001000100011010110100111010001" when "1010101011",
   "11010001011111010000111000010001011111111001000010110110011011001001100100" when "1010101100",
   "11010001011111010000111000010001011111111001000010110110011011001001100100" when "1010101101",
   "11010001101100100111000111011100101110000001011101110100110111110000111010" when "1010101110",
   "11010001111001111110000011001100101111001010101100010101100110110000100101" when "1010101111",
   "11010010000111010101101011100110001101010010100101101000110010000011011011" when "1010110000",
   "11010010000111010101101011100110001101010010100101101000110010000011011011" when "1010110001",
   "11010010010100101110000000101101110011000101101111000110111001010101011100" when "1010110010",
   "11010010100010000111000010101000001011111111100110000010011011001011011100" when "1010110011",
   "11010010100010000111000010101000001011111111100110000010011011001011011100" when "1010110100",
   "11010010101111100000110001011010000100001010101001011100000001111011101110" when "1010110101",
   "11010010111100111011001101001000001000100000100011111001010101001011011000" when "1010110110",
   "11010011001010010110010101110111000110101010010101011110010000100100000001" when "1010110111",
   "11010011001010010110010101110111000110101010010101011110010000100100000001" when "1010111000",
   "11010011010111110010001011101011101101000000011101101001000000110101110110" when "1010111001",
   "11010011100101001110101110101010101010101011000101010000100111111010101001" when "1010111010",
   "11010011100101001110101110101010101010101011000101010000100111111010101001" when "1010111011",
   "11010011110010101011111110111000101111100010001000100110001000101110010000" when "1010111100",
   "11010100000000001001111100011010101100001101100001011000011011110001100001" when "1010111101",
   "11010100000000001001111100011010101100001101100001011000011011110001100001" when "1010111110",
   "11010100001101101000100111010101010010000101010000111010101101001100111100" when "1010111111",
   "11010100011011000111111111101101010011010001101010001101100101001000110011" when "1011000000",
   "11010100101000101000000101100111100010101011011100001010111011010000100000" when "1011000001",
   "11010100101000101000000101100111100010101011011100001010111011010000100000" when "1011000010",
   "11010100110110001000111001001000110011111011111011110100010110010111010010" when "1011000011",
   "11010101000011101010011010010101111011011101001110100100011000110101000110" when "1011000100",
   "11010101000011101010011010010101111011011101001110100100011000110101000110" when "1011000101",
   "11010101010001001100101001010011101110011010010100100010011010110010001010" when "1011000110",
   "11010101011110101111100110000111000010101111010010111001010010111000100101" when "1011000111",
   "11010101011110101111100110000111000010101111010010111001010010111000100101" when "1011001000",
   "11010101101100010011010000110100101111001001011110010000101110100011100000" when "1011001001",
   "11010101111001110111101001100001101011000111100101001001011010100011010111" when "1011001010",
   "11010110000111011100110000010010101110111001111010011011111100101111101100" when "1011001011",
   "11010110000111011100110000010010101110111001111010011011111100101111101100" when "1011001100",
   "11010110010101000010100101001100110011100010011111111010011111111110101001" when "1011001101",
   "11010110100010101001001000010100110010110101010000110101010010111011010000" when "1011001110",
   "11010110100010101001001000010100110010110101010000110101010010111011010000" when "1011001111",
   "11010110110000010000011001101111100111011000001100100001111010110011010000" when "1011010000",
   "11010110111101111000011001100010001100100011100001000101011010110110001110" when "1011010001",
   "11010110111101111000011001100010001100100011100001000101011010110110001110" when "1011010010",
   "11010111001011100001000111110001011110100001110110000001010001011111100011" when "1011010011",
   "11010111011001001010100100100010011010010000010111000011001100000101100001" when "1011010100",
   "11010111011001001010100100100010011010010000010111000011001100000101100001" when "1011010101",
   "11010111100110110100101111111001111101011110111110110111110010000111110010" when "1011010110",
   "11010111110100011111101001111101000110110000100010000000001000111000010000" when "1011010111",
   "11010111110100011111101001111101000110110000100010000000001000111000010000" when "1011011000",
   "11011000000010001011010010110000110101011010111001101010010000011001010011" when "1011011001",
   "11011000001111110111101010011010001001100111001110101100011010101100111010" when "1011011010",
   "11011000011101100100110000111110000100010010000100100011011110010000100101" when "1011011011",
   "11011000011101100100110000111110000100010010000100100011011110010000100101" when "1011011100",
   "11011000101011010010100110100001100111001011100100010100000100100010000011" when "1011011101",
   "11011000111001000001001011001001110100110111100111101110110101101001100010" when "1011011110",
   "11011000111001000001001011001001110100110111100111101110110101101001100010" when "1011011111",
   "11011001000110110000011110111011110000101110000100010111100010000110010011" when "1011100000",
   "11011001010100100000100001111100011110111010110110101111001011011010110010" when "1011100001",
   "11011001010100100000100001111100011110111010110110101111001011011010110010" when "1011100010",
   "11011001100010010001010100010001000100011110001101100001001100110101110100" when "1011100011",
   "11011001110000000010110101111110100111001100110100110011100100110111001011" when "1011100100",
   "11011001110000000010110101111110100111001100110100110011100100110111001011" when "1011100101",
   "11011001111101110101000111001010001101110000000001011010000000101101011101" when "1011100110",
   "11011010001011101000000111111000111111100101111100001100001010101100001010" when "1011100111",
   "11011010001011101000000111111000111111100101111100001100001010101100001010" when "1011101000",
   "11011010011001011011111000010000000101000001101101011110111100011001000111" when "1011101001",
   "11011010100111010000011000010100100111001011101000100000110101110000011101" when "1011101010",
   "11011010100111010000011000010100100111001011101000100000110101110000011101" when "1011101011",
   "11011010110101000101101000001011110000000001010110111001011001111111010001" when "1011101100",
   "11011011000010111011100111111010101010010110000100001011110011010100110100" when "1011101101",
   "11011011000010111011100111111010101010010110000100001011110011010100110100" when "1011101110",
   "11011011010000110010010111100110100001110010101001011100011110101011000100" when "1011101111",
   "11011011011110101001110111010100100010110101111000111010000000000111100100" when "1011110000",
   "11011011011110101001110111010100100010110101111000111010000000000111100100" when "1011110001",
   "11011011101100100010000111001001111010110100101001101001000001010101110000" when "1011110010",
   "11011011111010011011000111001011110111111010000011010011011010111100101110" when "1011110011",
   "11011011111010011011000111001011110111111010000011010011011010111100101110" when "1011110100",
   "11011100001000010100110111011111101001000111101001111010101001110010010000" when "1011110101",
   "11011100010110001111011000001010011110010101101001101101010001001101111101" when "1011110110",
   "11011100010110001111011000001010011110010101101001101101010001001101111101" when "1011110111",
   "11011100100100001010101001010001101000010011000010111111101011011111010000" when "1011111000",
   "11011100110010000110101010111010011000100101110110001000001001001001011000" when "1011111001",
   "11011100110010000110101010111010011000100101110110001000001001001001011000" when "1011111010",
   "11011101000000000011011101001010000001101011001111011110000000101001011111" when "1011111011",
   "11011101001110000001000000000101110110110111110011011100001111001010100000" when "1011111100",
   "11011101001110000001000000000101110110110111110011011100001111001010100000" when "1011111101",
   "11011101011011111111010011110011001100010111101010100111001011101011110000" when "1011111110",
   "11011101101001111110011000010111010111001110101101110101101101011110110001" when "1011111111",
   "11011101101001111110011000010111010111001110101101110101101101011110110001" when "1100000000",
   "11011101110111111110001101110111101101011000110010011101100111000010000110" when "1100000001",
   "11011110000101111110110100011001100101101001110110100011010110011110100010" when "1100000010",
   "11011110000101111110110100011001100101101001110110100011010110011110100010" when "1100000011",
   "11011110010100000000001100000010010111101110001101001101001100101101000100" when "1100000100",
   "11011110010100000000001100000010010111101110001101001101001100101101000100" when "1100000101",
   "11011110100010000010010100110111011100001010101010111001101100001100001101" when "1100000110",
   "11011110110000000101001110111110001100011100110001111001100000101011100011" when "1100000111",
   "11011110110000000101001110111110001100011100110001111001100000101011100011" when "1100001000",
   "11011110111110001000111010011100000010111010111110101100110000110101001110" when "1100001001",
   "11011111001100001101010111010110011010110100110100100011101010111100111010" when "1100001010",
   "11011111001100001101010111010110011010110100110100100011101010111100111010" when "1100001011",
   "11011111011010010010100101110010110000010011001010000010101101111100110100" when "1100001100",
   "11011111101000011000100101110110100000011000010101101010001111101001011101" when "1100001101",
   "11011111101000011000100101110110100000011000010101101010001111101001011101" when "1100001110",
   "11011111110110011111010111100111001001000000011010100001100001100101001000" when "1100001111",
   "11100000000100100110111011001010001001000001010101000101010101011101000111" when "1100010000",
   "11100000000100100110111011001010001001000001010101000101010101011101000111" when "1100010001",
   "11100000010010101111010000100101000000001011000111111010000010011010010001" when "1100010010",
   "11100000010010101111010000100101000000001011000111111010000010011010010001" when "1100010011",
   "11100000100000111000010111111101001111001000001000100001001100001111110100" when "1100010100",
   "11100000101111000010010001011000010111011101001100010010101101110011001100" when "1100010101",
   "11100000101111000010010001011000010111011101001100010010101101110011001100" when "1100010110",
   "11100000111101001100111100111011111011101001110101011001100111101000001101" when "1100010111",
   "11100001001011011000011010101101011111001000011111110100010100001101110101" when "1100011000",
   "11100001001011011000011010101101011111001000011111110100010100001101110101" when "1100011001",
   "11100001011001100100101010110010100110001110101110011000100010110111011001" when "1100011010",
   "11100001100111110001101101010000110110001101010111111010111010011111011101" when "1100011011",
   "11100001100111110001101101010000110110001101010111111010111010011111011101" when "1100011100",
   "11100001110101111111100010001101110101010000110100011010000101100001010110" when "1100011101",
   "11100001110101111111100010001101110101010000110100011010000101100001010110" when "1100011110",
   "11100010000100001110001001101111001010100001001010001101101000000111001010" when "1100011111",
   "11100010010010011101100011111010011110000010011011011000100001111010100101" when "1100100000",
   "11100010010010011101100011111010011110000010011011011000100001111010100101" when "1100100001",
   "11100010100000101101110000110101011000110100110010111111011100100110111010" when "1100100010",
   "11100010101110111110110000100101100100110100110010100010101000011011110010" when "1100100011",
   "11100010101110111110110000100101100100110100110010100010101000011011110010" when "1100100100",
   "11100010111101010000100011010000101100111011011111011011101000000000000000" when "1100100101",
   "11100011001011100011001000111100011100111110110000011110101100100100101100" when "1100100110",
   "11100011001011100011001000111100011100111110110000011110101100100100101100" when "1100100111",
   "11100011011001110110100001101110100001110001011011100000000100001001011110" when "1100101000",
   "11100011011001110110100001101110100001110001011011100000000100001001011110" when "1100101001",
   "11100011101000001010101101101100101001000011100010111100111010100010101000" when "1100101010",
   "11100011110110011111101100111100100001100010100011101000001110110010111100" when "1100101011",
   "11100011110110011111101100111100100001100010100011101000001110110010111100" when "1100101100",
   "11100100000100110101011111100011111010111001100010011011011110001011011100" when "1100101101",
   "11100100010011001100000101101000100101110001011010001011000110000011010101" when "1100101110",
   "11100100010011001100000101101000100101110001011010001011000110000011010101" when "1100101111",
   "11100100100001100011011111010000010011110001001001011110111101111011110001" when "1100110000",
   "11100100100001100011011111010000010011110001001001011110111101111011110001" when "1100110001",
   "11100100101111111011101100100000110111011110000000101110101011000010011100" when "1100110010",
   "11100100111110010100101101100000000100011011110000000001101110100111110100" when "1100110011",
   "11100100111110010100101101100000000100011011110000000001101110100111110100" when "1100110100",
   "11100101001100101110100010010011101111001100110101010011110000011101000001" when "1100110101",
   "11100101001100101110100010010011101111001100110101010011110000011101000001" when "1100110110",
   "11100101011011001001001011000001101101010010101010011100100110101111010001" when "1100110111",
   "11100101101001100100100111101111110101001101110011011100011100110101110010" when "1100111000",
   "11100101101001100100100111101111110101001101110011011100011100110101110010" when "1100111001",
   "11100101111000000000111000100011111110011110001100101011111010001001001000" when "1100111010",
   "11100110000110011101111101100100000001100011011001010000001010011010010110" when "1100111011",
   "11100110000110011101111101100100000001100011011001010000001010011010010110" when "1100111100",
   "11100110010100111011110110110101110111111100110001010011001001000001001101" when "1100111101",
   "11100110010100111011110110110101110111111100110001010011001001000001001101" when "1100111110",
   "11100110100011011010100100011111011100001001110000011111110000011001101100" when "1100111111",
   "11100110110001111010000110100110101001101010000100100010001111001000110010" when "1101000000",
   "11100110110001111010000110100110101001101010000100100010001111001000110010" when "1101000001",
   "11100111000000011010011101010001011100111101111011101100100100000001101111" when "1101000010",
   "11100111000000011010011101010001011100111101111011101100100100000001101111" when "1101000011",
   "11100111001110111011101000100101110011100110010011011111000010100101001101" when "1101000100",
   "11100111011101011101101000101001101100000101000111010101000001010100010100" when "1101000101",
   "11100111011101011101101000101001101100000101000111010101000001010100010100" when "1101000110",
   "11100111101100000000011101100011000101111101011111010101110011010010010010" when "1101000111",
   "11100111101100000000011101100011000101111101011111010101110011010010010010" when "1101001000",
   "11100111111010100100000111011000000001110011111111001001101110001111110001" when "1101001001",
   "11101000001001001000100110001110100001001110110100110011011110111011101110" when "1101001010",
   "11101000001001001000100110001110100001001110110100110011011110111011101110" when "1101001011",
   "11101000010111101101111010001100100110110110000111101101101100110101111010" when "1101001100",
   "11101000010111101101111010001100100110110110000111101101101100110101111010" when "1101001101",
   "11101000100110010100000011011000010110010100000111101100101111000000001110" when "1101001110",
   "11101000110100111011000001110111110100010101011100000100110011001100000000" when "1101001111",
   "11101000110100111011000001110111110100010101011100000100110011001100000000" when "1101010000",
   "11101001000011100010110101110001000110101001010010110100011001000001101110" when "1101010001",
   "11101001000011100010110101110001000110101001010010110100011001000001101110" when "1101010010",
   "11101001010010001011011111001010010100000001101111110011000010100001001110" when "1101010011",
   "11101001100000110100111110001001100100010011111100000100011011011010010011" when "1101010100",
   "11101001100000110100111110001001100100010011111100000100011011011010010011" when "1101010101",
   "11101001101111011111010010110101000000011000010101001111111000111100111101" when "1101010110",
   "11101001101111011111010010110101000000011000010101001111111000111100111101" when "1101010111",
   "11101001111110001010011101010010110010001010111100111100010011100010000100" when "1101011000",
   "11101010001100110110011101101001000100101011101000010000011011101101011010" when "1101011001",
   "11101010001100110110011101101001000100101011101000010000011011101101011010" when "1101011010",
   "11101010011011100011010011111110000011111110001111010111101100001010100100" when "1101011011",
   "11101010011011100011010011111110000011111110001111010111101100001010100100" when "1101011100",
   "11101010101010010001000000010111111101001010111101001011011010000111001110" when "1101011101",
   "11101010111000111111100010111100111110011110011111000000100101101101100010" when "1101011110",
   "11101010111000111111100010111100111110011110011111000000100101101101100010" when "1101011111",
   "11101011000111101110111011110011010111001010010100011010001100000010000011" when "1101100000",
   "11101011000111101110111011110011010111001010010100011010001100000010000011" when "1101100001",
   "11101011010110011111001011000001010111100100111110111111111100001001100001" when "1101100010",
   "11101011010110011111001011000001010111100100111110111111111100001001100001" when "1101100011",
   "11101011100101010000010000101101010001001010010010011001110000111011000011" when "1101100100",
   "11101011110100000010001100111101010110011011100100001111110001000100010110" when "1101100101",
   "11101011110100000010001100111101010110011011100100001111110001000100010110" when "1101100110",
   "11101100000010110100111111110111111010111111111100001110110111000101101010" when "1101100111",
   "11101100000010110100111111110111111010111111111100001110110111000101101010" when "1101101000",
   "11101100010001101000101001100011010011100100100100010010000010101100101001" when "1101101001",
   "11101100100000011101001010000101110101111100111000110000010101010100110111" when "1101101010",
   "11101100100000011101001010000101110101111100111000110000010101010100110111" when "1101101011",
   "11101100101111010010100001100101111001000010111000101111011011010110011010" when "1101101100",
   "11101100101111010010100001100101111001000010111000101111011011010110011010" when "1101101101",
   "11101100111110001000110000001001110100110111010110011011000011101011000100" when "1101101110",
   "11101100111110001000110000001001110100110111010110011011000011101011000100" when "1101101111",
   "11101101001100111111110101111000000010100010000111100001000111010011010110" when "1101110000",
   "11101101011011110111110010110110111100010010010101110010100010100101011000" when "1101110001",
   "11101101011011110111110010110110111100010010010101110010100010100101011000" when "1101110010",
   "11101101101010110000100111001100111101011110101111101001000001110000010010" when "1101110011",
   "11101101101010110000100111001100111101011110101111101001000001110000010010" when "1101110100",
   "11101101111001101010010011000000100010100101111000110001100010011111100100" when "1101110101",
   "11101110001000100100110110011000001001001110011010111011101100001010000110" when "1101110110",
   "11101110001000100100110110011000001001001110011010111011101100001010000110" when "1101110111",
   "11101110010111100000010001011010010000000111010110101110000000011001111010" when "1101111000",
   "11101110010111100000010001011010010000000111010110101110000000011001111010" when "1101111001",
   "11101110100110011100100100001101010111001000010100011111000101111001110110" when "1101111010",
   "11101110100110011100100100001101010111001000010100011111000101111001110110" when "1101111011",
   "11101110110101011001101110110111111111010001110101010011101110110111010100" when "1101111100",
   "11101111000100010111110001100000101010101101100100000001111101000110110101" when "1101111101",
   "11101111000100010111110001100000101010101101100100000001111101000110110101" when "1101111110",
   "11101111010011010110101100001101111100101110100110011001000101011011000010" when "1101111111",
   "11101111010011010110101100001101111100101110100110011001000101011011000010" when "1110000000",
   "11101111100010010110011111000110011001110001101110001110110011111110010011" when "1110000001",
   "11101111100010010110011111000110011001110001101110001110110011111110010011" when "1110000010",
   "11101111110001010111001010010000100111011101101010110001010011011111110011" when "1110000011",
   "11110000000000011000101101110011001100100011011001111110011001000101111011" when "1110000100",
   "11110000000000011000101101110011001100100011011001111110011001000101111011" when "1110000101",
   "11110000001111011011001001110100110000111110011001111111110110011000001110" when "1110000110",
   "11110000001111011011001001110100110000111110011001111111110110011000001110" when "1110000111",
   "11110000011110011110011110011011111101110100111010101100110011110100000110" when "1110001000",
   "11110000011110011110011110011011111101110100111010101100110011110100000110" when "1110001001",
   "11110000101101100010101011101111011101011000001111010000010101000000001111" when "1110001010",
   "11110000101101100010101011101111011101011000001111010000010101000000001111" when "1110001011",
   "11110000111100100111110001110101111011000100111111110101001000110011001001" when "1110001100",
   "11110001001011101101110000110110000011100011011011010110100111000010011100" when "1110001101",
   "11110001001011101101110000110110000011100011011011010110100111000010011100" when "1110001110",
   "11110001011010110100101000110110100100100111101001010110111101110000111000" when "1110001111",
   "11110001011010110100101000110110100100100111101001010110111101110000111000" when "1110010000",
   "11110001101001111100011001111110001101010001111011111010101111110010000001" when "1110010001",
   "11110001101001111100011001111110001101010001111011111010101111110010000001" when "1110010010",
   "11110001111001000101000100010011101101101111000001101001100110011011001010" when "1110010011",
   "11110001111001000101000100010011101101101111000001101001100110011011001010" when "1110010100",
   "11110010001000001110100111111101110111011000010111110100011000011010010001" when "1110010101",
   "11110010010111011001000101000011011100110100011100100000100111101011100110" when "1110010110",
   "11110010010111011001000101000011011100110100011100100000100111101011100110" when "1110010111",
   "11110010100110100100011011101011010001110111000000111001011000001000100000" when "1110011000",
   "11110010100110100100011011101011010001110111000000111001011000001000100000" when "1110011001",
   "11110010110101110000101011111100001011100001011011100101100001001010000001" when "1110011010",
   "11110010110101110000101011111100001011100001011011100101100001001010000001" when "1110011011",
   "11110011000100111101110101111101000000000010111011000011011011111010110010" when "1110011100",
   "11110011000100111101110101111101000000000010111011000011011011111010110010" when "1110011101",
   "11110011010100001011111001110100100110111000111000001010010000010100110000" when "1110011110",
   "11110011100011011010110111101001111000101111001000110000100010100111111110" when "1110011111",
   "11110011100011011010110111101001111000101111001000110000100010100111111110" when "1110100000",
   "11110011110010101010101111100011101111100000010010011000100011101000010011" when "1110100001",
   "11110011110010101010101111100011101111100000010010011000100011101000010011" when "1110100010",
   "11110100000001111011100001101001000110010101111101000010000101100001000111" when "1110100011",
   "11110100000001111011100001101001000110010101111101000010000101100001000111" when "1110100100",
   "11110100010001001101001110000000111001101001000110000001110111001110010110" when "1110100101",
   "11110100010001001101001110000000111001101001000110000001110111001110010110" when "1110100110",
   "11110100100000011111110100110010000111000010010010111110101000011011111001" when "1110100111",
   "11110100101111110011010110000011101101011010000100110011111000001100000110" when "1110101000",
   "11110100101111110011010110000011101101011010000100110011111000001100000110" when "1110101001",
   "11110100111111000111110001111100101100111001001010111010010000001000000110" when "1110101010",
   "11110100111111000111110001111100101100111001001010111010010000001000000110" when "1110101011",
   "11110101001110011101001000100100000110111000110110010101101110011100101011" when "1110101100",
   "11110101001110011101001000100100000110111000110110010101101110011100101011" when "1110101101",
   "11110101011101110011011010000000111110000011001101001001100000100111101011" when "1110101110",
   "11110101011101110011011010000000111110000011001101001001100000100111101011" when "1110101111",
   "11110101101101001010100110011010010110010011011101110001110000111010110101" when "1110110000",
   "11110101101101001010100110011010010110010011011101110001110000111010110101" when "1110110001",
   "11110101111100100010101101110111010100110110010010100011001000111001100001" when "1110110010",
   "11110101111100100010101101110111010100110110010010100011001000111001100001" when "1110110011",
   "11110110001011111011110000011111000000001010000101010000001010110111111101" when "1110110100",
   "11110110011011010101101110011000011111111111010010110100100100100011011111" when "1110110101",
   "11110110011011010101101110011000011111111111010010110100100100100011011111" when "1110110110",
   "11110110101010110000100111101010111101011000101111000110011100111011110101" when "1110110111",
   "11110110101010110000100111101010111101011000101111000110011100111011110101" when "1110111000",
   "11110110111010001100011100011101100010101011111000101101011111100111000010" when "1110111001",
   "11110110111010001100011100011101100010101011111000101101011111100111000010" when "1110111010",
   "11110111001001101001001100110111011011100001001101000000000111101001101100" when "1110111011",
   "11110111001001101001001100110111011011100001001101000000000111101001101100" when "1110111100",
   "11110111011001000110111000111111110100110100011100000110101100001110110111" when "1110111101",
   "11110111011001000110111000111111110100110100011100000110101100001110110111" when "1110111110",
   "11110111101000100101100000111101111100110100111101000100110001001011011110" when "1110111111",
   "11110111101000100101100000111101111100110100111101000100110001001011011110" when "1111000000",
   "11110111111000000101000100111001000011000110000010001000011101101001111100" when "1111000001",
   "11111000000111100101100100111000011000011111001100111111111011001100000111" when "1111000010",
   "11111000000111100101100100111000011000011111001100111111111011001100000111" when "1111000011",
   "11111000010111000111000001000011001111001100100011010100111111010001111100" when "1111000100",
   "11111000010111000111000001000011001111001100100011010100111111010001111100" when "1111000101",
   "11111000100110101001011001100000111010101111000011001111000001110100110101" when "1111000110",
   "11111000100110101001011001100000111010101111000011001111000001110100110101" when "1111000111",
   "11111000110110001100101110011000101111111100110111111011000010101000001011" when "1111001000",
   "11111000110110001100101110011000101111111100110111111011000010101000001011" when "1111001001",
   "11111001000101110000111111110010000101000001101110011010000000010000101100" when "1111001010",
   "11111001000101110000111111110010000101000001101110011010000000010000101100" when "1111001011",
   "11111001010101010110001101110100010001011111001010010101100010100101000111" when "1111001100",
   "11111001010101010110001101110100010001011111001010010101100010100101000111" when "1111001101",
   "11111001100100111100011000100110101110001100111010111010111011001011111110" when "1111001110",
   "11111001100100111100011000100110101110001100111010111010111011001011111110" when "1111001111",
   "11111001110100100011100000010000110101011001001111111100011110001010100110" when "1111010000",
   "11111001110100100011100000010000110101011001001111111100011110001010100110" when "1111010001",
   "11111010000100001011100100111010000010101001001110111001010101011011011000" when "1111010010",
   "11111010000100001011100100111010000010101001001110111001010101011011011000" when "1111010011",
   "11111010010011110100100110101001110010111001001000001011110001000001011000" when "1111010100",
   "11111010100011011110100101100111100100011100101100011101110110110001000011" when "1111010101",
   "11111010100011011110100101100111100100011100101100011101110110110001000011" when "1111010110",
   "11111010110011001001100001111010110110111111100010000100110011100110100010" when "1111010111",
   "11111010110011001001100001111010110110111111100010000100110011100110100010" when "1111011000",
   "11111011000010110101011011101011001011100101011010100010110001000011001011" when "1111011001",
   "11111011000010110101011011101011001011100101011010100010110001000011001011" when "1111011010",
   "11111011010010100010010011000000000100101010101000001111010001001100110000" when "1111011011",
   "11111011010010100010010011000000000100101010101000001111010001001100110000" when "1111011100",
   "11111011100010010000001000000001000110000100010100000110010011101010000100" when "1111011101",
   "11111011100010010000001000000001000110000100010100000110010011101010000100" when "1111011110",
   "11111011110001111110111010110101110101000000110011011110000101111001110000" when "1111011111",
   "11111011110001111110111010110101110101000000110011011110000101111001110000" when "1111100000",
   "11111100000001101110101011100101111000000111111110000011100001100000110001" when "1111100001",
   "11111100000001101110101011100101111000000111111110000011100001100000110001" when "1111100010",
   "11111100010001011111011010011000110111011011100011111101011010101111100010" when "1111100011",
   "11111100010001011111011010011000110111011011100011111101011010101111100010" when "1111100100",
   "11111100100001010001000111010110011100010111100011110110100001111101101000" when "1111100101",
   "11111100100001010001000111010110011100010111100011110110100001111101101000" when "1111100110",
   "11111100110001000011110010100110010001110010100001001110011010011100110110" when "1111100111",
   "11111100110001000011110010100110010001110010100001001110011010011100110110" when "1111101000",
   "11111101000000110111011100010000000011111101111010110001001001000101101101" when "1111101001",
   "11111101000000110111011100010000000011111101111010110001001001000101101101" when "1111101010",
   "11111101010000101100000100011011100000100110100000110101111101100000101010" when "1111101011",
   "11111101010000101100000100011011100000100110100000110101111101100000101010" when "1111101100",
   "11111101100000100001101011010000010110110100101100000100111000001111111110" when "1111101101",
   "11111101100000100001101011010000010110110100101100000100111000001111111110" when "1111101110",
   "11111101110000011000010000110110010111001100110100000011010000011111111111" when "1111101111",
   "11111101110000011000010000110110010111001100110100000011010000011111111111" when "1111110000",
   "11111110000000001111110101010101010011101111100110000111011100000011110010" when "1111110001",
   "11111110000000001111110101010101010011101111100110000111011100000011110010" when "1111110010",
   "11111110010000001000011000110100111111111010011100010011011100000110010110" when "1111110011",
   "11111110010000001000011000110100111111111010011100010011011100000110010110" when "1111110100",
   "11111110100000000001111011011101010000100111110100010110110001011000011111" when "1111110101",
   "11111110100000000001111011011101010000100111110100010110110001011000011111" when "1111110110",
   "11111110101111111100011101010101111100001111100110110111011010100101101100" when "1111110111",
   "11111110101111111100011101010101111100001111100110110111011010100101101100" when "1111111000",
   "11111110111111110111111110100110111010100111011110100001111111011010111111" when "1111111001",
   "11111110111111110111111110100110111010100111011110100001111111011010111111" when "1111111010",
   "11111111001111110100011111011000000101000011001111100001001011001011101100" when "1111111011",
   "11111111001111110100011111011000000101000011001111100001001011001011101100" when "1111111100",
   "11111111011111110001111111110001010110010101001110111100011001100001110110" when "1111111101",
   "11111111011111110001111111110001010110010101001110111100011001100001110110" when "1111111110",
   "11111111101111110000011111111010101010101110101010011101111000001000100000" when "1111111111",
   "--------------------------------------------------------------------------" when others;
    Y <= TableOut_d1;
end architecture;

--------------------------------------------------------------------------------
--                         LogTable_1_8_66_F400_uid76
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity LogTable_1_8_66_F400_uid76 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          Y : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of LogTable_1_8_66_F400_uid76 is
signal TableOut :  std_logic_vector(65 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "000000001000000000000000000111111111111111110101010101010101100101" when "00000000",
   "000000011000000000000000001000000000000000001010101010101010111011" when "00000001",
   "000000101000000000000001001000000000000100100000000000010100010000" when "00000010",
   "000000111000000000000011001000000000010100110101010111110001100110" when "00000011",
   "000001001000000000000110001000000000111001001010110100000010111100" when "00000100",
   "000001011000000000001010001000000001111001100000011001101000010110" when "00000101",
   "000001101000000000001111001000000011011101110110001110100001110101" when "00000110",
   "000001111000000000010101001000000101101110001100011010001111011111" when "00000111",
   "000010001000000000011100001000001000110010100011000101110001011010" when "00001000",
   "000010011000000000100100001000001100110010111010011011100111110000" when "00001001",
   "000010101000000000101101001000010001110111010010100111110010101100" when "00001010",
   "000010111000000000110111001000011000000111101011110111110010011111" when "00001011",
   "000011001000000001000010001000011111101100000110011010100111011010" when "00001100",
   "000011011000000001001110001000101000101100100010100000110001110100" when "00001101",
   "000011101000000001011011001000110011010001000000011100010010001010" when "00001110",
   "000011111000000001101001001000111111100001100000100000101000111001" when "00001111",
   "000100001000000001111000001001001101100110000011000010110110100111" when "00010000",
   "000100011000000010001000001001011101100110101000011001011011111111" when "00010001",
   "000100101000000010011001001001101111101011010000111100011001110000" when "00010010",
   "000100111000000010101011001010000011111011111101000101010000110000" when "00010011",
   "000101001000000010111110001010011010100000101101001111000001111101" when "00010100",
   "000101011000000011010010001010110011100001100001110110001110011010" when "00010101",
   "000101101000000011100111001011001111000110011011011000110111010011" when "00010110",
   "000101111000000011111101001011101101010111011010010110011101111010" when "00010111",
   "000110001000000100010100001100001110011100011111010000000011101001" when "00011000",
   "000110011000000100101100001100110010011101101010101000001010000101" when "00011001",
   "000110101000000101000101001101011001100010111101000010110010111001" when "00011010",
   "000110111000000101011111001110000011110100010111000101011111111010" when "00011011",
   "000111001000000101111010001110110001011001111001010111010011001001" when "00011100",
   "000111011000000110010110001111100010011011100100100000101110101100" when "00011101",
   "000111101000000110110011010000010111000001011001001011110100111000" when "00011110",
   "000111111000000111010001010001001111010011011000000100001000001011" when "00011111",
   "001000001000000111110000010010001011011001100001110110101011001100" when "00100000",
   "001000011000001000010000010011001011011011110111010010000000110010" when "00100001",
   "001000101000001000110001010100001111100010011001000110001011111011" when "00100010",
   "001000111000001001010011010101010111110101001000000100101111110100" when "00100011",
   "001001001000001001110110010110100100011100000101000000101111110111" when "00100100",
   "001001011000001010011010010111110101011111010000101110101111101001" when "00100101",
   "001001101000001010111111011001001011000110101100000100110010111110" when "00100110",
   "001001111000001011100101011010100101011010010111111010011101110101" when "00100111",
   "001010001000001100001100011100000100100010010101001000110100100000" when "00101000",
   "001010011000001100110100011101101000100110100100101010011011011010" when "00101001",
   "001010101000001101011101011111010001101111000111011011010111010000" when "00101010",
   "001010111000001110000111100001000000000011111110011001001100111111" when "00101011",
   "001011001000001110110010100010110011101101001010100011000001110000" when "00101100",
   "001011011000001111011110100100101100110010101100111001011011000000" when "00101101",
   "001011101000010000001011100110101011011100100110011110011110011010" when "00101110",
   "001011111000010000111001101000101111110010111000010101110001111001" when "00101111",
   "001100001000010001101000101010111001111101100011100100011011101100" when "00110000",
   "001100011000010010011000101101001010000100101001010001000010010000" when "00110001",
   "001100101000010011001001101111100000010000001010100011101100010110" when "00110010",
   "001100111000010011111011110001111100101000001000100110000001000010" when "00110011",
   "001101001000010100101110110100011111010100100100100011000111101000" when "00110100",
   "001101011000010101100010110111001000011101011111100111100111110001" when "00110101",
   "001101101000010110010111111001111000001010111011000001101001011001" when "00110110",
   "001101111000010111001101111100101110100100111000000000110100101111" when "00110111",
   "001110001000011000000100111111101011110011010111110110010010010111" when "00111000",
   "001110011000011000111101000010101111111110011011110100101011001000" when "00111001",
   "001110101000011001110110000101111011001110000101010000001000010000" when "00111010",
   "001110111000011010110000001001001101101010010101011110010011010000" when "00111011",
   "001111001000011011101011001100100111011011001101110110010110000001" when "00111100",
   "001111011000011100100111010000001000101000101111110000111010110000" when "00111101",
   "001111101000011101100100010011110001011010111100101000001100000010" when "00111110",
   "001111111000011110100010010111100001111001110101110111110100110000" when "00111111",
   "010000001000011111100001011011011010001101011100111101000000001101" when "01000000",
   "010000011000100000100001011111011010011101110011010110011010000011" when "01000001",
   "010000101000100001100010100011100010110010111010100100001110010010" when "01000010",
   "010000111000100010100100100111110011010100110100001000001001010100" when "01000011",
   "010001001000100011100111101100001100001011100001100101010111111100" when "01000100",
   "010001011000100100101011110000101101011111000100100000100111010101" when "01000101",
   "010001101000100101110000110101010111010111011110100000000101000011" when "01000110",
   "010001111000100110110110111010001001111100110001001011011111000100" when "01000111",
   "010010001000100111111101111111000101010110111110001100000011110001" when "01001000",
   "010010011000101001000110000100001001101110000111001100100001111100" when "01001001",
   "010010101000101010001111001001010111001010001101111001001000110101" when "01001010",
   "010010111000101011011001001110101101110011010011111111101000000011" when "01001011",
   "010011001000101100100100010100001101110001011011001111001111101100" when "01001100",
   "010011011000101101110000011001110111001100100101011000110000010000" when "01001101",
   "010011101000101110111101011111101010001100110100001110011010101100" when "01001110",
   "010011111000110000001011100101100110111010001001100100000000011010" when "01001111",
   "010100001000110001011010101011101101011100100111001110110011010010" when "01010000",
   "010100011000110010101010110001111101111100001111000101100101101000" when "01010001",
   "010100101000110011111011111000011000100001000011000000101010001110" when "01010010",
   "010100111000110101001101111110111101010011000100111001110100010100" when "01010011",
   "010101001000110110100001000101101100011010010110101100010111101100" when "01010100",
   "010101011000110111110101001100100101111110111010010101001000100100" when "01010101",
   "010101101000111001001010010011101010001000110001110010011011101000" when "01010110",
   "010101111000111010100000011010111000111111111111000100000110000110" when "01010111",
   "010110001000111011110111100010010010101100100100001011011101101101" when "01011000",
   "010110011000111101001111101001110111010110100011001011011000101010" when "01011001",
   "010110101000111110101000110001100111000101111110001000001101101111" when "01011010",
   "010110111001000000000010111001100010000010110111000111110100001010" when "01011011",
   "010111001001000001011110000001101000010101010000010001100011101110" when "01011100",
   "010111011001000010111010001001111010000101001011101110010100101110" when "01011101",
   "010111101001000100010111010010010111011010101011101000100000000100" when "01011110",
   "010111111001000101110101011011000000011101110010001011111111000111" when "01011111",
   "011000001001000111010100100011110101010110100001100110001011110100" when "01100000",
   "011000011001001000110100101100110110001100111100000110000000101101" when "01100001",
   "011000101001001010010101110110000011001001000011111011111000110100" when "01100010",
   "011000111001001011110111111111011100010010111011011001101111110100" when "01100011",
   "011001001001001101011011001001000001110010100100110011000001111000" when "01100100",
   "011001011001001110111111010010110011110000000010011100101011110011" when "01100101",
   "011001101001010000100100011100110010010011010110101101001010111110" when "01100110",
   "011001111001010010001010100110111101100100100011111100011101010110" when "01100111",
   "011010001001010011110001110001010101101011101100100100000001011110" when "01101000",
   "011010011001010101011001111011111010110000110010111110110110100001" when "01101001",
   "011010101001010111000011000110101100111011111001101001011100010001" when "01101010",
   "011010111001011000101101010001101100010101000011000001110011000110" when "01101011",
   "011011001001011010011000011100111001000100010001100111011100000010" when "01101100",
   "011011011001011100000100101000010011010001100111111011011000101011" when "01101101",
   "011011101001011101110001110011111011000101001000100000001011010100" when "01101110",
   "011011111001011111011111111111110000100110110101111001110110110111" when "01101111",
   "011100001001100001001111001011110011111110110010101101111110110110" when "01110000",
   "011100011001100010111111011000000101010101000001100011100111011110" when "01110001",
   "011100101001100100110000100100100100110001100101000011010101100111" when "01110010",
   "011100111001100110100010110001010010011100011111110111001110110001" when "01110011",
   "011101001001101000010101111110001110011101110100101010111001001000" when "01110100",
   "011101011001101010001010001011011000111101100110001011011011100100" when "01110101",
   "011101101001101011111111011000110010000011110111000111011101100110" when "01110110",
   "011101111001101101110101100110011001111000101010001111000111011100" when "01110111",
   "011110001001101111101100110100010000100100000010010100000010000011" when "01111000",
   "011110011001110001100101000010010110001110000010001001010111000001" when "01111001",
   "011110101001110011011110010000101010111110101100100011110000101010" when "01111010",
   "011110111001110101011000011111001110111110000100011001011010000000" when "01111011",
   "011111001001110111010011101110000010010100001100100001111110110010" when "01111100",
   "011111011001111001001111111101000101001001000111110110101011011111" when "01111101",
   "011111101001111011001101001100010111100100111001010010001101010010" when "01111110",
   "011111111001111101001011011011111001101111100011110000110010000110" when "01111111",
   "100000000001111110001010111011110000110000111111010100011100011100" when "10000000",
   "100000010010000000001010101011101010110001000100111011110011100001" when "10000001",
   "100000100010000010001011011011110100110100001011000011010111101010" when "10000010",
   "100000110010000100001101001100001111000010010100101100101001011011" when "10000011",
   "100001000010000110001111111100111001100011100100111010101010000101" when "10000100",
   "100001010010001000010011101101110100011111111110110001111011101101" when "10000101",
   "100001100010001010011000011110111111111111100101011000100001001000" when "10000110",
   "100001110010001100011110010000011100001010011011110101111101111101" when "10000111",
   "100010000010001110100101000010001001001000100101010011010110100101" when "10001000",
   "100010010010010000101100110100000111000010000100111011010000001011" when "10001001",
   "100010100010010010110101100110010101111110111101111001110000101111" when "10001010",
   "100010110010010100111111011000110110000111010011011100011111000001" when "10001011",
   "100011000010010111001010001011100111100011001000110010100010101000" when "10001100",
   "100011010010011001010101111110101010011010100001001100100011111100" when "10001101",
   "100011100010011011100010110001111110110101011111111100101100001100" when "10001110",
   "100011110010011101110000100101100100111100001000010110100101011010" when "10001111",
   "100100000010011111111111011001011100110110011101101111011010011111" when "10010000",
   "100100010010100010001111001101100110101100100011011101110111000110" when "10010001",
   "100100100010100100100000000010000010100110011100111010000111110011" when "10010010",
   "100100110010100110110001110110110000101100001101011101111010000001" when "10010011",
   "100101000010101001000100101011110001000101111000100100011011111111" when "10010100",
   "100101010010101011011000100001000011111011100001101010011100110100" when "10010101",
   "100101100010101101101101010110101001010101001100001110001100100000" when "10010110",
   "100101110010110000000011001100100001011010111011101111011011111000" when "10010111",
   "100110000010110010011010000010101100010100110011101111011100101100" when "10011000",
   "100110010010110100110001111001001010001010110111110001000001100010" when "10011001",
   "100110100010110111001010101111111011000101001011011000011101111011" when "10011010",
   "100110110010111001100100100110111111001011110010001011100110010000" when "10011011",
   "100111000010111011111111011110010110100110101111110001101111110110" when "10011100",
   "100111010010111110011011010110000001011110000111110011110000111000" when "10011101",
   "100111100011000000111000001101111111111001111101111100000000011111" when "10011110",
   "100111110011000011010110000110010010000010010101110110010110101110" when "10011111",
   "101000000011000101110100111110110111111111010011010000001100100011" when "10100000",
   "101000010011001000010100110111110001111000111001111000011011110110" when "10100001",
   "101000100011001010110101110000111111110111001101011111011111011110" when "10100010",
   "101000110011001101010111101010100010000010010001110111010011001101" when "10100011",
   "101001000011001111111010100100011000100010001010110011010011110000" when "10100100",
   "101001010011010010011110011110100011011110111100001000011110110101" when "10100101",
   "101001100011010101000011011001000011000000101001101101010011000011" when "10100110",
   "101001110011010111101001010011110111001111010111011001110000000011" when "10100111",
   "101010000011011010010000001111000000010011001001000111010110011010" when "10101000",
   "101010010011011100111000001010011110010100000010110001000111101011" when "10101001",
   "101010100011011111100001000110010001011010001000010011100110011010" when "10101010",
   "101010110011100010001011000010011001101101011101101100110110001001" when "10101011",
   "101011000011100100110101111110110111010110000110111100011011011011" when "10101100",
   "101011010011100111100001111011101010011100001000000011011011110010" when "10101101",
   "101011100011101010001110111000110011000111100101000100011101110010" when "10101110",
   "101011110011101100111100110110010001100000100010000011101000111101" when "10101111",
   "101100000011101111101011110100000101101111000011000110100101111001" when "10110000",
   "101100010011110010011011110010001111111011001100010100011110001101" when "10110001",
   "101100100011110101001100110000110000001101000001110101111100100011" when "10110010",
   "101100110011110111111110101111100110101100100111110101001100100100" when "10110011",
   "101101000011111010110001101110110011100010000010011101111011000001" when "10110100",
   "101101010011111101100101101110010110110101010101111101010101101010" when "10110101",
   "101101100100000000011010101110010000101110100110100010001011010100" when "10110110",
   "101101110100000011010000101110100001010101111000011100101011111000" when "10110111",
   "101110000100000110000111101111001000110011001111111110101000010100" when "10111000",
   "101110010100001000111111110000000111001110110001011011010010101001" when "10111001",
   "101110100100001011111000110001011100110000100001000111011101111111" when "10111010",
   "101110110100001110110010110011001001100000100011011001011110100011" when "10111011",
   "101111000100010001101101110101001101100110111100101001001001100111" when "10111100",
   "101111010100010100101001110111101001001011110001001111110101100011" when "10111101",
   "101111100100010111100110111010011100010111000101101000011001111000" when "10111110",
   "101111110100011010100100111101100111010000111110001111001111001100" when "10111111",
   "110000000100011101100100000001001010000001011111100010001111001011" when "11000000",
   "110000010100100000100100000101000100110000101110000000110100101101" when "11000001",
   "110000100100100011100101001001010111100110101110001011111011101111" when "11000010",
   "110000110100100110100111001110000010101011100100100110000001010111" when "11000011",
   "110001000100101001101010010011000110000111010101110011000011110011" when "11000100",
   "110001010100101100101110011000100010000010000110011000100010011110" when "11000101",
   "110001100100101111110011011110010110100011111010111101011101111000" when "11000110",
   "110001110100110010111001100100100011110100111000001010010111101111" when "11000111",
   "110010000100110110000000101011001001111101000010101001010010110111" when "11001000",
   "110010010100111001001000110010001001000100011111000101110011010100" when "11001001",
   "110010100100111100010001111001100001010011010010001100111110010010" when "11001010",
   "110010110100111111011100000001010010110001100000101101011010001000" when "11001011",
   "110011000101000010100111001001011101100111001111010111001110011100" when "11001100",
   "110011010101000101110011010010000001111100100010111100000011111101" when "11001101",
   "110011100101001001000000011010111111111001100000001111000100101000" when "11001110",
   "110011110101001100001110100100010111100110001100000100111011101001" when "11001111",
   "110100000101001111011101101110001001001010101011010011110101010111" when "11010000",
   "110100010101010010101101111000010100101111000010110011011111010111" when "11010001",
   "110100100101010101111111000010111010011011010111011101001000011101" when "11010010",
   "110100110101011001010001001101111010010111101110001011100000101101" when "11010011",
   "110101000101011100100100011001010100101100001011111010111001010111" when "11010100",
   "110101010101011111111000100101001001100000110101101001000100111100" when "11010101",
   "110101100101100011001101110001011000111101110000010101010111001101" when "11010110",
   "110101110101100110100011111110000011001011000001000000100101001011" when "11010111",
   "110110000101101001111011001011001000010000101100101101000101001000" when "11011000",
   "110110010101101101010011011000101000010110111000011110101110100101" when "11011001",
   "110110100101110000101100100110100011100101101001011010111010010110" when "11011010",
   "110110110101110100000110110100111010000101000100101000100010100000" when "11011011",
   "110111000101110111100010000011101011111101001111010000000010011011" when "11011100",
   "110111010101111010111110010010111001010110001110011011010110110000" when "11011101",
   "110111100101111110011011100010100010011000000111010101111101011011" when "11011110",
   "110111110110000001111001110010100111001010111111001100110101101110" when "11011111",
   "111000000110000101011001000011000111110110111011001110100000001010" when "11100000",
   "111000010110001000111001010100000100100100000000101010111110100111" when "11100001",
   "111000100110001100011010100101011101011010010100110011110100010001" when "11100010",
   "111000110110001111111100110111010010100001111100111100000101100111" when "11100011",
   "111001000110010011100000001001100100000010111110011000011000100001" when "11100100",
   "111001010110010111000100011100010010000101011110011110110100000111" when "11100101",
   "111001100110011010101001101111011100110001100010100111000000111100" when "11100110",
   "111001110110011110010000000011000100001111010000001010001000110110" when "11100111",
   "111010000110100001110111010111001000100110101100100010110111000010" when "11101000",
   "111010010110100101011111101011101001111111111101001101011000000110" when "11101001",
   "111010100110101001001001000000101000100011000111100111011001111110" when "11101010",
   "111010110110101100110011010110000100011000010001010000001011111101" when "11101011",
   "111011000110110000011110101011111101100111011111101000011110110000" when "11101100",
   "111011010110110100001011000010010100011000111000010010100100011010" when "11101101",
   "111011100110110111111000011001001000110100100000110010010000011010" when "11101110",
   "111011110110111011100110110000011011000010011110101100110111100110" when "11101111",
   "111100000110111111010110001000001011001010110111101001010000001111" when "11110000",
   "111100010111000011000110100000011001010101110001001111110001111111" when "11110001",
   "111100100111000110110111111001000101101011010001001010010101111011" when "11110010",
   "111100110111001010101010010010010000010011011101000100010110100011" when "11110011",
   "111101000111001110011101101011111001010110011010101010101111110010" when "11110100",
   "111101010111010010010010000110000000111100001111101011111110111110" when "11110101",
   "111101100111010110000111100000100111001101000001111000000010111010" when "11110110",
   "111101110111011001111101111011101100010000110111000000011011110110" when "11110111",
   "111110000111011101110101010111010000001111110100111000001011011100" when "11111000",
   "111110010111100001101101110011010011010010000001010011110100110101" when "11111001",
   "111110100111100101100111001111110101011111100010001001011100101000" when "11111010",
   "111110110111101001100001101100110111000000011101010000101000111010" when "11111011",
   "111111000111101101011101001010010111111100111000100010100001001011" when "11111100",
   "111111010111110001011001101000011000011100111001111001101110011110" when "11111101",
   "111111100111110101010111000110111000101000100111010010011011010011" when "11111110",
   "111111110111111001010101100101111000101000000110101010010011101001" when "11111111",
   "------------------------------------------------------------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_74_f400_uid80
--                    (IntAdderAlternative_74_F400_uid84)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_74_f400_uid80 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(73 downto 0);
          Y : in  std_logic_vector(73 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(73 downto 0)   );
end entity;

architecture arch of IntAdder_74_f400_uid80 is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(32 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(31 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(32 downto 0);
signal sum_l1_idx1 :  std_logic_vector(31 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(73 downto 42)) + ( "0" & Y(73 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
   sum_l0_idx1 <= s_sum_l0_idx1(31 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(32 downto 32);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(31 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(32 downto 32);
   R <= sum_l1_idx1(31 downto 0) & sum_l0_idx0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        LogTable_2_10_59_F400_uid88
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity LogTable_2_10_59_F400_uid88 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(58 downto 0)   );
end entity;

architecture arch of LogTable_2_10_59_F400_uid88 is
signal TableOut :  std_logic_vector(58 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "00000000000000000000000000000000000000000000010000000000000" when "0000000000",
   "00000000010000000000000000000000000011110000010000000000000" when "0000000001",
   "00000000100000000000000000000000001111100000010000000000001" when "0000000010",
   "00000000110000000000000000000000100011010000010000000000100" when "0000000011",
   "00000001000000000000000000000000111111000000010000000001010" when "0000000100",
   "00000001010000000000000000000001100010110000010000000010100" when "0000000101",
   "00000001100000000000000000000010001110100000010000000100011" when "0000000110",
   "00000001110000000000000000000011000010010000010000000111000" when "0000000111",
   "00000010000000000000000000000011111110000000010000001010100" when "0000001000",
   "00000010010000000000000000000101000001110000010000001111000" when "0000001001",
   "00000010100000000000000000000110001101100000010000010100101" when "0000001010",
   "00000010110000000000000000000111100001010000010000011011100" when "0000001011",
   "00000011000000000000000000001000111101000000010000100011110" when "0000001100",
   "00000011010000000000000000001010100000110000010000101101100" when "0000001101",
   "00000011100000000000000000001100001100100000010000111000110" when "0000001110",
   "00000011110000000000000000001110000000010000010001000101111" when "0000001111",
   "00000100000000000000000000001111111100000000010001010100111" when "0000010000",
   "00000100010000000000000000010001111111110000010001100101110" when "0000010001",
   "00000100100000000000000000010100001011100000010001111000111" when "0000010010",
   "00000100110000000000000000010110011111010000010010001110010" when "0000010011",
   "00000101000000000000000000011000111011000000010010100101111" when "0000010100",
   "00000101010000000000000000011011011110110000010011000000001" when "0000010101",
   "00000101100000000000000000011110001010100000010011011100111" when "0000010110",
   "00000101110000000000000000100000111110010000010011111100100" when "0000010111",
   "00000110000000000000000000100011111010000000010100011110111" when "0000011000",
   "00000110010000000000000000100110111101110000010101000100010" when "0000011001",
   "00000110100000000000000000101010001001100000010101101100111" when "0000011010",
   "00000110110000000000000000101101011101010000010110011000101" when "0000011011",
   "00000111000000000000000000110000111001000000010111000111110" when "0000011100",
   "00000111010000000000000000110100011100110000010111111010100" when "0000011101",
   "00000111100000000000000000111000001000100000011000110000110" when "0000011110",
   "00000111110000000000000000111011111100010000011001101010110" when "0000011111",
   "00001000000000000000000000111111111000000000011010101000101" when "0000100000",
   "00001000010000000000000001000011111011110000011011101010100" when "0000100001",
   "00001000100000000000000001001000000111100000011100110000101" when "0000100010",
   "00001000110000000000000001001100011011010000011101111010111" when "0000100011",
   "00001001000000000000000001010000110111000000011111001001100" when "0000100100",
   "00001001010000000000000001010101011010110000100000011100101" when "0000100101",
   "00001001100000000000000001011010000110100000100001110100011" when "0000100110",
   "00001001110000000000000001011110111010010000100011010000111" when "0000100111",
   "00001010000000000000000001100011110110000000100100110010010" when "0000101000",
   "00001010010000000000000001101000111001110000100110011000101" when "0000101001",
   "00001010100000000000000001101110000101100000101000000100000" when "0000101010",
   "00001010110000000000000001110011011001010000101001110100110" when "0000101011",
   "00001011000000000000000001111000110101000000101011101010111" when "0000101100",
   "00001011010000000000000001111110011000110000101101100110100" when "0000101101",
   "00001011100000000000000010000100000100100000101111100111110" when "0000101110",
   "00001011110000000000000010001001111000010000110001101110101" when "0000101111",
   "00001100000000000000000010001111110100000000110011111011100" when "0000110000",
   "00001100010000000000000010010101110111110000110110001110011" when "0000110001",
   "00001100100000000000000010011100000011100000111000100111010" when "0000110010",
   "00001100110000000000000010100010010111010000111011000110100" when "0000110011",
   "00001101000000000000000010101000110011000000111101101100000" when "0000110100",
   "00001101010000000000000010101111010110110001000000011000001" when "0000110101",
   "00001101100000000000000010110110000010100001000011001010110" when "0000110110",
   "00001101110000000000000010111100110110010001000110000100010" when "0000110111",
   "00001110000000000000000011000011110010000001001001000100100" when "0000111000",
   "00001110010000000000000011001010110101110001001100001011111" when "0000111001",
   "00001110100000000000000011010010000001100001001111011010010" when "0000111010",
   "00001110110000000000000011011001010101010001010010110000000" when "0000111011",
   "00001111000000000000000011100000110001000001010110001101000" when "0000111100",
   "00001111010000000000000011101000010100110001011001110001100" when "0000111101",
   "00001111100000000000000011110000000000100001011101011101101" when "0000111110",
   "00001111110000000000000011110111110100010001100001010001101" when "0000111111",
   "00010000000000000000000011111111110000000001100101001101011" when "0001000000",
   "00010000010000000000000100000111110011110001101001010001001" when "0001000001",
   "00010000100000000000000100001111111111100001101101011101000" when "0001000010",
   "00010000110000000000000100011000010011010001110001110001001" when "0001000011",
   "00010001000000000000000100100000101111000001110110001101101" when "0001000100",
   "00010001010000000000000100101001010010110001111010110010101" when "0001000101",
   "00010001100000000000000100110001111110100001111111100000010" when "0001000110",
   "00010001110000000000000100111010110010010010000100010110101" when "0001000111",
   "00010010000000000000000101000011101110000010001001010101111" when "0001001000",
   "00010010010000000000000101001100110001110010001110011110001" when "0001001001",
   "00010010100000000000000101010101111101100010010011101111100" when "0001001010",
   "00010010110000000000000101011111010001010010011001001010001" when "0001001011",
   "00010011000000000000000101101000101101000010011110101110001" when "0001001100",
   "00010011010000000000000101110010010000110010100100011011100" when "0001001101",
   "00010011100000000000000101111011111100100010101010010010101" when "0001001110",
   "00010011110000000000000110000101110000010010110000010011100" when "0001001111",
   "00010100000000000000000110001111101100000010110110011110010" when "0001010000",
   "00010100010000000000000110011001101111110010111100110010111" when "0001010001",
   "00010100100000000000000110100011111011100011000011010001110" when "0001010010",
   "00010100110000000000000110101110001111010011001001111010110" when "0001010011",
   "00010101000000000000000110111000101011000011010000101110010" when "0001010100",
   "00010101010000000000000111000011001110110011010111101100010" when "0001010101",
   "00010101100000000000000111001101111010100011011110110100110" when "0001010110",
   "00010101110000000000000111011000101110010011100110001000000" when "0001010111",
   "00010110000000000000000111100011101010000011101101100110010" when "0001011000",
   "00010110010000000000000111101110101101110011110101001111011" when "0001011001",
   "00010110100000000000000111111001111001100011111101000011110" when "0001011010",
   "00010110110000000000001000000101001101010100000101000011010" when "0001011011",
   "00010111000000000000001000010000101001000100001101001110001" when "0001011100",
   "00010111010000000000001000011100001100110100010101100100101" when "0001011101",
   "00010111100000000000001000100111111000100100011110000110101" when "0001011110",
   "00010111110000000000001000110011101100010100100110110100011" when "0001011111",
   "00011000000000000000001000111111101000000100101111101110000" when "0001100000",
   "00011000010000000000001001001011101011110100111000110011110" when "0001100001",
   "00011000100000000000001001010111110111100101000010000101100" when "0001100010",
   "00011000110000000000001001100100001011010101001011100011100" when "0001100011",
   "00011001000000000000001001110000100111000101010101001101111" when "0001100100",
   "00011001010000000000001001111101001010110101011111000100110" when "0001100101",
   "00011001100000000000001010001001110110100101101001001000010" when "0001100110",
   "00011001110000000000001010010110101010010101110011011000100" when "0001100111",
   "00011010000000000000001010100011100110000101111101110101101" when "0001101000",
   "00011010010000000000001010110000101001110110001000011111110" when "0001101001",
   "00011010100000000000001010111101110101100110010011010111000" when "0001101010",
   "00011010110000000000001011001011001001010110011110011011100" when "0001101011",
   "00011011000000000000001011011000100101000110101001101101010" when "0001101100",
   "00011011010000000000001011100110001000110110110101001100101" when "0001101101",
   "00011011100000000000001011110011110100100111000000111001101" when "0001101110",
   "00011011110000000000001100000001101000010111001100110100011" when "0001101111",
   "00011100000000000000001100001111100100000111011000111100111" when "0001110000",
   "00011100010000000000001100011101100111110111100101010011100" when "0001110001",
   "00011100100000000000001100101011110011100111110001111000010" when "0001110010",
   "00011100110000000000001100111010000111010111111110101011001" when "0001110011",
   "00011101000000000000001101001000100011001000001011101100100" when "0001110100",
   "00011101010000000000001101010111000110111000011000111100010" when "0001110101",
   "00011101100000000000001101100101110010101000100110011010110" when "0001110110",
   "00011101110000000000001101110100100110011000110100000111111" when "0001110111",
   "00011110000000000000001110000011100010001001000010000100000" when "0001111000",
   "00011110010000000000001110010010100101111001010000001111000" when "0001111001",
   "00011110100000000000001110100001110001101001011110101001010" when "0001111010",
   "00011110110000000000001110110001000101011001101101010010101" when "0001111011",
   "00011111000000000000001111000000100001001001111100001011011" when "0001111100",
   "00011111010000000000001111010000000100111010001011010011110" when "0001111101",
   "00011111100000000000001111011111110000101010011010101011101" when "0001111110",
   "00011111110000000000001111101111100100011010101010010011010" when "0001111111",
   "00100000000000000000001111111111100000001010111010001010110" when "0010000000",
   "00100000010000000000010000001111100011111011001010010010010" when "0010000001",
   "00100000100000000000010000011111101111101011011010101010000" when "0010000010",
   "00100000110000000000010000110000000011011011101011010001111" when "0010000011",
   "00100001000000000000010001000000011111001011111100001010001" when "0010000100",
   "00100001010000000000010001010001000010111100001101010010111" when "0010000101",
   "00100001100000000000010001100001101110101100011110101100010" when "0010000110",
   "00100001110000000000010001110010100010011100110000010110011" when "0010000111",
   "00100010000000000000010010000011011110001101000010010001011" when "0010001000",
   "00100010010000000000010010010100100001111101010100011101011" when "0010001001",
   "00100010100000000000010010100101101101101101100110111010100" when "0010001010",
   "00100010110000000000010010110111000001011101111001101000111" when "0010001011",
   "00100011000000000000010011001000011101001110001100101000100" when "0010001100",
   "00100011010000000000010011011010000000111110011111111001110" when "0010001101",
   "00100011100000000000010011101011101100101110110011011100101" when "0010001110",
   "00100011110000000000010011111101100000011111000111010001010" when "0010001111",
   "00100100000000000000010100001111011100001111011011010111110" when "0010010000",
   "00100100010000000000010100100001011111111111101111110000001" when "0010010001",
   "00100100100000000000010100110011101011110000000100011010110" when "0010010010",
   "00100100110000000000010101000101111111100000011001010111101" when "0010010011",
   "00100101000000000000010101011000011011010000101110100110110" when "0010010100",
   "00100101010000000000010101101010111111000001000100001000100" when "0010010101",
   "00100101100000000000010101111101101010110001011001111100110" when "0010010110",
   "00100101110000000000010110010000011110100001110000000011111" when "0010010111",
   "00100110000000000000010110100011011010010010000110011101110" when "0010011000",
   "00100110010000000000010110110110011110000010011101001010110" when "0010011001",
   "00100110100000000000010111001001101001110010110100001010110" when "0010011010",
   "00100110110000000000010111011100111101100011001011011110001" when "0010011011",
   "00100111000000000000010111110000011001010011100011000100110" when "0010011100",
   "00100111010000000000011000000011111101000011111010111110111" when "0010011101",
   "00100111100000000000011000010111101000110100010011001100110" when "0010011110",
   "00100111110000000000011000101011011100100100101011101110010" when "0010011111",
   "00101000000000000000011000111111011000010101000100100011101" when "0010100000",
   "00101000010000000000011001010011011100000101011101101101000" when "0010100001",
   "00101000100000000000011001100111100111110101110111001010100" when "0010100010",
   "00101000110000000000011001111011111011100110010000111100011" when "0010100011",
   "00101001000000000000011010010000010111010110101011000010100" when "0010100100",
   "00101001010000000000011010100100111011000111000101011101001" when "0010100101",
   "00101001100000000000011010111001100110110111100000001100011" when "0010100110",
   "00101001110000000000011011001110011010100111111011010000011" when "0010100111",
   "00101010000000000000011011100011010110011000010110101001010" when "0010101000",
   "00101010010000000000011011111000011010001000110010010111001" when "0010101001",
   "00101010100000000000011100001101100101111001001110011010001" when "0010101010",
   "00101010110000000000011100100010111001101001101010110010011" when "0010101011",
   "00101011000000000000011100111000010101011010000111100000000" when "0010101100",
   "00101011010000000000011101001101111001001010100100100011000" when "0010101101",
   "00101011100000000000011101100011100100111011000001111011110" when "0010101110",
   "00101011110000000000011101111001011000101011011111101010010" when "0010101111",
   "00101100000000000000011110001111010100011011111101101110101" when "0010110000",
   "00101100010000000000011110100101011000001100011100001001000" when "0010110001",
   "00101100100000000000011110111011100011111100111010111001100" when "0010110010",
   "00101100110000000000011111010001110111101101011010000000001" when "0010110011",
   "00101101000000000000011111101000010011011101111001011101010" when "0010110100",
   "00101101010000000000011111111110110111001110011001010000110" when "0010110101",
   "00101101100000000000100000010101100010111110111001011011000" when "0010110110",
   "00101101110000000000100000101100010110101111011001111100000" when "0010110111",
   "00101110000000000000100001000011010010011111111010110011110" when "0010111000",
   "00101110010000000000100001011010010110010000011100000010100" when "0010111001",
   "00101110100000000000100001110001100010000000111101101000100" when "0010111010",
   "00101110110000000000100010001000110101110001011111100101110" when "0010111011",
   "00101111000000000000100010100000010001100010000001111010010" when "0010111100",
   "00101111010000000000100010110111110101010010100100100110010" when "0010111101",
   "00101111100000000000100011001111100001000011000111101010000" when "0010111110",
   "00101111110000000000100011100111010100110011101011000101011" when "0010111111",
   "00110000000000000000100011111111010000100100001110111000101" when "0011000000",
   "00110000010000000000100100010111010100010100110011000100000" when "0011000001",
   "00110000100000000000100100101111100000000101010111100111011" when "0011000010",
   "00110000110000000000100101000111110011110101111100100011000" when "0011000011",
   "00110001000000000000100101100000001111100110100001110111000" when "0011000100",
   "00110001010000000000100101111000110011010111000111100011100" when "0011000101",
   "00110001100000000000100110010001011111000111101101101000101" when "0011000110",
   "00110001110000000000100110101010010010111000010100000110100" when "0011000111",
   "00110010000000000000100111000011001110101000111010111101010" when "0011001000",
   "00110010010000000000100111011100010010011001100010001101000" when "0011001001",
   "00110010100000000000100111110101011110001010001001110110000" when "0011001010",
   "00110010110000000000101000001110110001111010110001111000000" when "0011001011",
   "00110011000000000000101000101000001101101011011010010011100" when "0011001100",
   "00110011010000000000101001000001110001011100000011001000100" when "0011001101",
   "00110011100000000000101001011011011101001100101100010111001" when "0011001110",
   "00110011110000000000101001110101010000111101010101111111100" when "0011001111",
   "00110100000000000000101010001111001100101110000000000001110" when "0011010000",
   "00110100010000000000101010101001010000011110101010011110000" when "0011010001",
   "00110100100000000000101011000011011100001111010101010100010" when "0011010010",
   "00110100110000000000101011011101110000000000000000100100111" when "0011010011",
   "00110101000000000000101011111000001011110000101100001111111" when "0011010100",
   "00110101010000000000101100010010101111100001011000010101010" when "0011010101",
   "00110101100000000000101100101101011011010010000100110101011" when "0011010110",
   "00110101110000000000101101001000001111000010110001110000010" when "0011010111",
   "00110110000000000000101101100011001010110011011111000101111" when "0011011000",
   "00110110010000000000101101111110001110100100001100110110101" when "0011011001",
   "00110110100000000000101110011001011010010100111011000010011" when "0011011010",
   "00110110110000000000101110110100101110000101101001101001100" when "0011011011",
   "00110111000000000000101111010000001001110110011000101011111" when "0011011100",
   "00110111010000000000101111101011101101100111001000001001111" when "0011011101",
   "00110111100000000000110000000111011001010111111000000011011" when "0011011110",
   "00110111110000000000110000100011001101001000101000011000110" when "0011011111",
   "00111000000000000000110000111111001000111001011001001001111" when "0011100000",
   "00111000010000000000110001011011001100101010001010010111000" when "0011100001",
   "00111000100000000000110001110111011000011010111100000000010" when "0011100010",
   "00111000110000000000110010010011101100001011101110000101111" when "0011100011",
   "00111001000000000000110010110000000111111100100000100111110" when "0011100100",
   "00111001010000000000110011001100101011101101010011100110001" when "0011100101",
   "00111001100000000000110011101001010111011110000111000001001" when "0011100110",
   "00111001110000000000110100000110001011001110111010111001000" when "0011100111",
   "00111010000000000000110100100011000110111111101111001101100" when "0011101000",
   "00111010010000000000110101000000001010110000100011111111010" when "0011101001",
   "00111010100000000000110101011101010110100001011001001110000" when "0011101010",
   "00111010110000000000110101111010101010010010001110111010000" when "0011101011",
   "00111011000000000000110110011000000110000011000101000011011" when "0011101100",
   "00111011010000000000110110110101101001110011111011101010010" when "0011101101",
   "00111011100000000000110111010011010101100100110010101110110" when "0011101110",
   "00111011110000000000110111110001001001010101101010010001000" when "0011101111",
   "00111100000000000000111000001111000101000110100010010001000" when "0011110000",
   "00111100010000000000111000101101001000110111011010101111001" when "0011110001",
   "00111100100000000000111001001011010100101000010011101011011" when "0011110010",
   "00111100110000000000111001101001101000011001001101000101111" when "0011110011",
   "00111101000000000000111010001000000100001010000110111110110" when "0011110100",
   "00111101010000000000111010100110100111111011000001010110000" when "0011110101",
   "00111101100000000000111011000101010011101011111100001100000" when "0011110110",
   "00111101110000000000111011100100000111011100110111100000110" when "0011110111",
   "00111110000000000000111100000011000011001101110011010100010" when "0011111000",
   "00111110010000000000111100100010000110111110101111100110111" when "0011111001",
   "00111110100000000000111101000001010010101111101100011000101" when "0011111010",
   "00111110110000000000111101100000100110100000101001101001100" when "0011111011",
   "00111111000000000000111110000000000010010001100111011001111" when "0011111100",
   "00111111010000000000111110011111100110000010100101101001110" when "0011111101",
   "00111111100000000000111110111111010001110011100100011001001" when "0011111110",
   "00111111110000000000111111011111000101100100100011101000010" when "0011111111",
   "01000000000000000000111111111111000001010101100011010111011" when "0100000000",
   "01000000010000000001000000011111000101000110100011100110011" when "0100000001",
   "01000000100000000001000000111111010000110111100100010101100" when "0100000010",
   "01000000110000000001000001011111100100101000100101100101000" when "0100000011",
   "01000001000000000001000010000000000000011001100111010100110" when "0100000100",
   "01000001010000000001000010100000100100001010101001100101000" when "0100000101",
   "01000001100000000001000011000001001111111011101100010110000" when "0100000110",
   "01000001110000000001000011100010000011101100101111100111101" when "0100000111",
   "01000010000000000001000100000010111111011101110011011010001" when "0100001000",
   "01000010010000000001000100100100000011001110110111101101110" when "0100001001",
   "01000010100000000001000101000101001110111111111100100010010" when "0100001010",
   "01000010110000000001000101100110100010110001000001111000010" when "0100001011",
   "01000011000000000001000110000111111110100010000111101111100" when "0100001100",
   "01000011010000000001000110101001100010010011001110001000010" when "0100001101",
   "01000011100000000001000111001011001110000100010101000010101" when "0100001110",
   "01000011110000000001000111101101000001110101011100011110110" when "0100001111",
   "01000100000000000001001000001110111101100110100100011100110" when "0100010000",
   "01000100010000000001001000110001000001010111101100111100110" when "0100010001",
   "01000100100000000001001001010011001101001000110101111110110" when "0100010010",
   "01000100110000000001001001110101100000111001111111100011010" when "0100010011",
   "01000101000000000001001010010111111100101011001001101010000" when "0100010100",
   "01000101010000000001001010111010100000011100010100010011010" when "0100010101",
   "01000101100000000001001011011101001100001101011111011111000" when "0100010110",
   "01000101110000000001001011111111111111111110101011001101101" when "0100010111",
   "01000110000000000001001100100010111011101111110111011111000" when "0100011000",
   "01000110010000000001001101000101111111100001000100010011100" when "0100011001",
   "01000110100000000001001101101001001011010010010001101011001" when "0100011010",
   "01000110110000000001001110001100011111000011011111100110000" when "0100011011",
   "01000111000000000001001110101111111010110100101110000100010" when "0100011100",
   "01000111010000000001001111010011011110100101111101000101111" when "0100011101",
   "01000111100000000001001111110111001010010111001100101011010" when "0100011110",
   "01000111110000000001010000011010111110001000011100110100010" when "0100011111",
   "01001000000000000001010000111110111001111001101101100001010" when "0100100000",
   "01001000010000000001010001100010111101101010111110110010010" when "0100100001",
   "01001000100000000001010010000111001001011100010000100111010" when "0100100010",
   "01001000110000000001010010101011011101001101100011000000100" when "0100100011",
   "01001001000000000001010011001111111000111110110101111110010" when "0100100100",
   "01001001010000000001010011110100011100110000001001100000011" when "0100100101",
   "01001001100000000001010100011001001000100001011101100111010" when "0100100110",
   "01001001110000000001010100111101111100010010110010010010110" when "0100100111",
   "01001010000000000001010101100010111000000100000111100011001" when "0100101000",
   "01001010010000000001010110000111111011110101011101011000100" when "0100101001",
   "01001010100000000001010110101101000111100110110011110011000" when "0100101010",
   "01001010110000000001010111010010011011011000001010110010111" when "0100101011",
   "01001011000000000001010111110111110111001001100010011000000" when "0100101100",
   "01001011010000000001011000011101011010111010111010100010101" when "0100101101",
   "01001011100000000001011001000011000110101100010011010011000" when "0100101110",
   "01001011110000000001011001101000111010011101101100101001000" when "0100101111",
   "01001100000000000001011010001110110110001111000110100100110" when "0100110000",
   "01001100010000000001011010110100111010000000100001000110110" when "0100110001",
   "01001100100000000001011011011011000101110001111100001110110" when "0100110010",
   "01001100110000000001011100000001011001100011010111111101000" when "0100110011",
   "01001101000000000001011100100111110101010100110100010001100" when "0100110100",
   "01001101010000000001011101001110011001000110010001001100110" when "0100110101",
   "01001101100000000001011101110101000100110111101110101110100" when "0100110110",
   "01001101110000000001011110011011111000101001001100110111000" when "0100110111",
   "01001110000000000001011111000010110100011010101011100110010" when "0100111000",
   "01001110010000000001011111101001111000001100001010111100110" when "0100111001",
   "01001110100000000001100000010001000011111101101010111010001" when "0100111010",
   "01001110110000000001100000111000010111101111001011011110111" when "0100111011",
   "01001111000000000001100001011111110011100000101100101011000" when "0100111100",
   "01001111010000000001100010000111010111010010001110011110100" when "0100111101",
   "01001111100000000001100010101111000011000011110000111001110" when "0100111110",
   "01001111110000000001100011010110110110110101010011111100110" when "0100111111",
   "01010000000000000001100011111110110010100110110111100111100" when "0101000000",
   "01010000010000000001100100100110110110011000011011111010011" when "0101000001",
   "01010000100000000001100101001111000010001010000000110101011" when "0101000010",
   "01010000110000000001100101110111010101111011100110011000100" when "0101000011",
   "01010001000000000001100110011111110001101101001100100100001" when "0101000100",
   "01010001010000000001100111001000010101011110110011011000010" when "0101000101",
   "01010001100000000001100111110001000001010000011010110100111" when "0101000110",
   "01010001110000000001101000011001110101000010000010111010010" when "0101000111",
   "01010010000000000001101001000010110000110011101011101000101" when "0101001000",
   "01010010010000000001101001101011110100100101010101000000000" when "0101001001",
   "01010010100000000001101010010101000000010110111111000000011" when "0101001010",
   "01010010110000000001101010111110010100001000101001101010000" when "0101001011",
   "01010011000000000001101011100111101111111010010100111101000" when "0101001100",
   "01010011010000000001101100010001010011101100000000111001101" when "0101001101",
   "01010011100000000001101100111010111111011101101101011111110" when "0101001110",
   "01010011110000000001101101100100110011001111011010101111110" when "0101001111",
   "01010100000000000001101110001110101111000001001000101001100" when "0101010000",
   "01010100010000000001101110111000110010110010110111001101010" when "0101010001",
   "01010100100000000001101111100010111110100100100110011011001" when "0101010010",
   "01010100110000000001110000001101010010010110010110010011010" when "0101010011",
   "01010101000000000001110000110111101110001000000110110101110" when "0101010100",
   "01010101010000000001110001100010010001111001111000000010110" when "0101010101",
   "01010101100000000001110010001100111101101011101001111010100" when "0101010110",
   "01010101110000000001110010110111110001011101011100011100110" when "0101010111",
   "01010110000000000001110011100010101101001111001111101010000" when "0101011000",
   "01010110010000000001110100001101110001000001000011100010010" when "0101011001",
   "01010110100000000001110100111000111100110010111000000101110" when "0101011010",
   "01010110110000000001110101100100010000100100101101010100010" when "0101011011",
   "01010111000000000001110110001111101100010110100011001110010" when "0101011100",
   "01010111010000000001110110111011010000001000011001110011110" when "0101011101",
   "01010111100000000001110111100110111011111010010001000101000" when "0101011110",
   "01010111110000000001111000010010101111101100001001000001110" when "0101011111",
   "01011000000000000001111000111110101011011110000001101010100" when "0101100000",
   "01011000010000000001111001101010101111001111111010111111010" when "0101100001",
   "01011000100000000001111010010110111011000001110101000000000" when "0101100010",
   "01011000110000000001111011000011001110110011101111101101010" when "0101100011",
   "01011001000000000001111011101111101010100101101011000110101" when "0101100100",
   "01011001010000000001111100011100001110010111100111001100101" when "0101100101",
   "01011001100000000001111101001000111010001001100011111111010" when "0101100110",
   "01011001110000000001111101110101101101111011100001011110100" when "0101100111",
   "01011010000000000001111110100010101001101101011111101010110" when "0101101000",
   "01011010010000000001111111001111101101011111011110100100000" when "0101101001",
   "01011010100000000001111111111100111001010001011110001010010" when "0101101010",
   "01011010110000000010000000101010001101000011011110011101110" when "0101101011",
   "01011011000000000010000001010111101000110101011111011110110" when "0101101100",
   "01011011010000000010000010000101001100100111100001001101010" when "0101101101",
   "01011011100000000010000010110010111000011001100011101001010" when "0101101110",
   "01011011110000000010000011100000101100001011100110110011000" when "0101101111",
   "01011100000000000010000100001110100111111101101010101010110" when "0101110000",
   "01011100010000000010000100111100101011101111101111010000011" when "0101110001",
   "01011100100000000010000101101010110111100001110100100100010" when "0101110010",
   "01011100110000000010000110011001001011010011111010100110010" when "0101110011",
   "01011101000000000010000111000111100111000110000001010110101" when "0101110100",
   "01011101010000000010000111110110001010111000001000110101100" when "0101110101",
   "01011101100000000010001000100100110110101010010001000011001" when "0101110110",
   "01011101110000000010001001010011101010011100011001111111011" when "0101110111",
   "01011110000000000010001010000010100110001110100011101010100" when "0101111000",
   "01011110010000000010001010110001101010000000101110000100110" when "0101111001",
   "01011110100000000010001011100000110101110010111001001110000" when "0101111010",
   "01011110110000000010001100010000001001100101000101000110100" when "0101111011",
   "01011111000000000010001100111111100101010111010001101110011" when "0101111100",
   "01011111010000000010001101101111001001001001011111000101110" when "0101111101",
   "01011111100000000010001110011110110100111011101101001100110" when "0101111110",
   "01011111110000000010001111001110101000101101111100000011100" when "0101111111",
   "01100000000000000010001111111110100100100000001011101010001" when "0110000000",
   "01100000010000000010010000101110101000010010011100000000110" when "0110000001",
   "01100000100000000010010001011110110100000100101101000111100" when "0110000010",
   "01100000110000000010010010001111000111110110111110111110100" when "0110000011",
   "01100001000000000010010010111111100011101001010001100101111" when "0110000100",
   "01100001010000000010010011110000000111011011100100111101110" when "0110000101",
   "01100001100000000010010100100000110011001101111001000110010" when "0110000110",
   "01100001110000000010010101010001100111000000001101111111100" when "0110000111",
   "01100010000000000010010110000010100010110010100011101001100" when "0110001000",
   "01100010010000000010010110110011100110100100111010000100110" when "0110001001",
   "01100010100000000010010111100100110010010111010001010000111" when "0110001010",
   "01100010110000000010011000010110000110001001101001001110011" when "0110001011",
   "01100011000000000010011001000111100001111100000001111101010" when "0110001100",
   "01100011010000000010011001111001000101101110011011011101100" when "0110001101",
   "01100011100000000010011010101010110001100000110101101111100" when "0110001110",
   "01100011110000000010011011011100100101010011010000110011010" when "0110001111",
   "01100100000000000010011100001110100001000101101100101000110" when "0110010000",
   "01100100010000000010011101000000100100111000001001010000011" when "0110010001",
   "01100100100000000010011101110010110000101010100110101010000" when "0110010010",
   "01100100110000000010011110100101000100011101000100110110000" when "0110010011",
   "01100101000000000010011111010111100000001111100011110100010" when "0110010100",
   "01100101010000000010100000001010000100000010000011100101001" when "0110010101",
   "01100101100000000010100000111100101111110100100100001000100" when "0110010110",
   "01100101110000000010100001101111100011100111000101011110110" when "0110010111",
   "01100110000000000010100010100010011111011001100111100111110" when "0110011000",
   "01100110010000000010100011010101100011001100001010100011111" when "0110011001",
   "01100110100000000010100100001000101110111110101110010011000" when "0110011010",
   "01100110110000000010100100111100000010110001010010110101100" when "0110011011",
   "01100111000000000010100101101111011110100011111000001011010" when "0110011100",
   "01100111010000000010100110100011000010010110011110010100100" when "0110011101",
   "01100111100000000010100111010110101110001001000101010001100" when "0110011110",
   "01100111110000000010101000001010100001111011101101000010001" when "0110011111",
   "01101000000000000010101000111110011101101110010101100110101" when "0110100000",
   "01101000010000000010101001110010100001100000111110111111010" when "0110100001",
   "01101000100000000010101010100110101101010011101001001011110" when "0110100010",
   "01101000110000000010101011011011000001000110010100001100110" when "0110100011",
   "01101001000000000010101100001111011100111001000000000010000" when "0110100100",
   "01101001010000000010101101000100000000101011101100101011110" when "0110100101",
   "01101001100000000010101101111000101100011110011010001010001" when "0110100110",
   "01101001110000000010101110101101100000010001001000011101010" when "0110100111",
   "01101010000000000010101111100010011100000011110111100101010" when "0110101000",
   "01101010010000000010110000010111011111110110100111100010010" when "0110101001",
   "01101010100000000010110001001100101011101001011000010100100" when "0110101010",
   "01101010110000000010110010000001111111011100001001111011110" when "0110101011",
   "01101011000000000010110010110111011011001110111100011000100" when "0110101100",
   "01101011010000000010110011101100111111000001101111101010110" when "0110101101",
   "01101011100000000010110100100010101010110100100011110010101" when "0110101110",
   "01101011110000000010110101011000011110100111011000110000010" when "0110101111",
   "01101100000000000010110110001110011010011010001110100011110" when "0110110000",
   "01101100010000000010110111000100011110001101000101001101010" when "0110110001",
   "01101100100000000010110111111010101001111111111100101100110" when "0110110010",
   "01101100110000000010111000110000111101110010110101000010110" when "0110110011",
   "01101101000000000010111001100111011001100101101110001110111" when "0110110100",
   "01101101010000000010111010011101111101011000101000010001101" when "0110110101",
   "01101101100000000010111011010100101001001011100011001011000" when "0110110110",
   "01101101110000000010111100001011011100111110011110111011000" when "0110110111",
   "01101110000000000010111101000010011000110001011011100010000" when "0110111000",
   "01101110010000000010111101111001011100100100011001000000000" when "0110111001",
   "01101110100000000010111110110000101000010111010111010101000" when "0110111010",
   "01101110110000000010111111100111111100001010010110100001011" when "0110111011",
   "01101111000000000011000000011111010111111101010110100101000" when "0110111100",
   "01101111010000000011000001010110111011110000010111100000010" when "0110111101",
   "01101111100000000011000010001110100111100011011001010011001" when "0110111110",
   "01101111110000000011000011000110011011010110011011111101110" when "0110111111",
   "01110000000000000011000011111110010111001001011111100000001" when "0111000000",
   "01110000010000000011000100110110011010111100100011111010100" when "0111000001",
   "01110000100000000011000101101110100110101111101001001101001" when "0111000010",
   "01110000110000000011000110100110111010100010101111011000000" when "0111000011",
   "01110001000000000011000111011111010110010101110110011011001" when "0111000100",
   "01110001010000000011001000010111111010001000111110010110110" when "0111000101",
   "01110001100000000011001001010000100101111100000111001011000" when "0111000110",
   "01110001110000000011001010001001011001101111010000111000001" when "0111000111",
   "01110010000000000011001011000010010101100010011011011110000" when "0111001000",
   "01110010010000000011001011111011011001010101100110111101000" when "0111001001",
   "01110010100000000011001100110100100101001000110011010101000" when "0111001010",
   "01110010110000000011001101101101111000111100000000100110010" when "0111001011",
   "01110011000000000011001110100111010100101111001110110001000" when "0111001100",
   "01110011010000000011001111100000111000100010011101110101000" when "0111001101",
   "01110011100000000011010000011010100100010101101101110010111" when "0111001110",
   "01110011110000000011010001010100011000001000111110101010011" when "0111001111",
   "01110100000000000011010010001110010011111100010000011011110" when "0111010000",
   "01110100010000000011010011001000010111101111100011000111010" when "0111010001",
   "01110100100000000011010100000010100011100010110110101100110" when "0111010010",
   "01110100110000000011010100111100110111010110001011001100100" when "0111010011",
   "01110101000000000011010101110111010011001001100000100110100" when "0111010100",
   "01110101010000000011010110110001110110111100110110111011010" when "0111010101",
   "01110101100000000011010111101100100010110000001110001010100" when "0111010110",
   "01110101110000000011011000100111010110100011100110010100100" when "0111010111",
   "01110110000000000011011001100010010010010110111111011001010" when "0111011000",
   "01110110010000000011011010011101010110001010011001011001010" when "0111011001",
   "01110110100000000011011011011000100001111101110100010100010" when "0111011010",
   "01110110110000000011011100010011110101110001010000001010100" when "0111011011",
   "01110111000000000011011101001111010001100100101100111100000" when "0111011100",
   "01110111010000000011011110001010110101011000001010101001010" when "0111011101",
   "01110111100000000011011111000110100001001011101001010010000" when "0111011110",
   "01110111110000000011100000000010010100111111001000110110011" when "0111011111",
   "01111000000000000011100000111110010000110010101001010110110" when "0111100000",
   "01111000010000000011100001111010010100100110001010110011000" when "0111100001",
   "01111000100000000011100010110110100000011001101101001011100" when "0111100010",
   "01111000110000000011100011110010110100001101010000100000010" when "0111100011",
   "01111001000000000011100100101111010000000000110100110001011" when "0111100100",
   "01111001010000000011100101101011110011110100011001111111000" when "0111100101",
   "01111001100000000011100110101000011111101000000000001001010" when "0111100110",
   "01111001110000000011100111100101010011011011100111010000001" when "0111100111",
   "01111010000000000011101000100010001111001111001111010100000" when "0111101000",
   "01111010010000000011101001011111010011000010111000010100110" when "0111101001",
   "01111010100000000011101010011100011110110110100010010010110" when "0111101010",
   "01111010110000000011101011011001110010101010001101001110000" when "0111101011",
   "01111011000000000011101100010111001110011101111001000110100" when "0111101100",
   "01111011010000000011101101010100110010010001100101111100101" when "0111101101",
   "01111011100000000011101110010010011110000101010011110000010" when "0111101110",
   "01111011110000000011101111010000010001111001000010100001110" when "0111101111",
   "01111100000000000011110000001110001101101100110010010001000" when "0111110000",
   "01111100010000000011110001001100010001100000100010111110011" when "0111110001",
   "01111100100000000011110010001010011101010100010100101001110" when "0111110010",
   "01111100110000000011110011001000110001001000000111010011100" when "0111110011",
   "01111101000000000011110100000111001100111011111010111011100" when "0111110100",
   "01111101010000000011110101000101110000101111101111100010000" when "0111110101",
   "01111101100000000011110110000100011100100011100101000111010" when "0111110110",
   "01111101110000000011110111000011010000010111011011101011001" when "0111110111",
   "01111110000000000011111000000010001100001011010011001110000" when "0111111000",
   "01111110010000000011111001000001001111111111001011101111110" when "0111111001",
   "01111110100000000011111010000000011011110011000101010000101" when "0111111010",
   "01111110110000000011111010111111101111100110111111110000110" when "0111111011",
   "01111111000000000011111011111111001011011010111011010000010" when "0111111100",
   "01111111010000000011111100111110101111001110110111101111011" when "0111111101",
   "01111111100000000011111101111110011011000010110101001110000" when "0111111110",
   "01111111110000000011111110111110001110110110110011101100100" when "0111111111",
   "10000000000000000011111111111110001010101010110011001010110" when "1000000000",
   "10000000010000000100000000111110001110011110110011101001000" when "1000000001",
   "10000000100000000100000001111110011010010010110101000111011" when "1000000010",
   "10000000110000000100000010111110101110000110110111100110000" when "1000000011",
   "10000001000000000100000011111111001001111010111011000101000" when "1000000100",
   "10000001010000000100000100111111101101101110111111100100100" when "1000000101",
   "10000001100000000100000110000000011001100011000101000100101" when "1000000110",
   "10000001110000000100000111000001001101010111001011100101100" when "1000000111",
   "10000010000000000100001000000010001001001011010011000111010" when "1000001000",
   "10000010010000000100001001000011001100111111011011101010000" when "1000001001",
   "10000010100000000100001010000100011000110011100101001101111" when "1000001010",
   "10000010110000000100001011000101101100100111101111110011000" when "1000001011",
   "10000011000000000100001100000111001000011011111011011001100" when "1000001100",
   "10000011010000000100001101001000101100010000001000000001100" when "1000001101",
   "10000011100000000100001110001010011000000100010101101011001" when "1000001110",
   "10000011110000000100001111001100001011111000100100010110100" when "1000001111",
   "10000100000000000100010000001110000111101100110100000011110" when "1000010000",
   "10000100010000000100010001010000001011100001000100110011000" when "1000010001",
   "10000100100000000100010010010010010111010101010110100100010" when "1000010010",
   "10000100110000000100010011010100101011001001101001010111111" when "1000010011",
   "10000101000000000100010100010111000110111101111101001101111" when "1000010100",
   "10000101010000000100010101011001101010110010010010000110011" when "1000010101",
   "10000101100000000100010110011100010110100110101000000001100" when "1000010110",
   "10000101110000000100010111011111001010011010111110111111010" when "1000010111",
   "10000110000000000100011000100010000110001111010111000000000" when "1000011000",
   "10000110010000000100011001100101001010000011110000000011110" when "1000011001",
   "10000110100000000100011010101000010101111000001010001010100" when "1000011010",
   "10000110110000000100011011101011101001101100100101010100101" when "1000011011",
   "10000111000000000100011100101111000101100001000001100010001" when "1000011100",
   "10000111010000000100011101110010101001010101011110110011000" when "1000011101",
   "10000111100000000100011110110110010101001001111101000111101" when "1000011110",
   "10000111110000000100011111111010001000111110011100100000000" when "1000011111",
   "10001000000000000100100000111110000100110010111100111100001" when "1000100000",
   "10001000010000000100100010000010001000100111011110011100011" when "1000100001",
   "10001000100000000100100011000110010100011100000001000000101" when "1000100010",
   "10001000110000000100100100001010101000010000100100101001010" when "1000100011",
   "10001001000000000100100101001111000100000101001001010110001" when "1000100100",
   "10001001010000000100100110010011100111111001101111000111101" when "1000100101",
   "10001001100000000100100111011000010011101110010101111101101" when "1000100110",
   "10001001110000000100101000011101000111100010111101111000100" when "1000100111",
   "10001010000000000100101001100010000011010111100110111000001" when "1000101000",
   "10001010010000000100101010100111000111001100010000111100110" when "1000101001",
   "10001010100000000100101011101100010011000000111100000110101" when "1000101010",
   "10001010110000000100101100110001100110110101101000010101101" when "1000101011",
   "10001011000000000100101101110111000010101010010101101010001" when "1000101100",
   "10001011010000000100101110111100100110011111000100000100000" when "1000101101",
   "10001011100000000100110000000010010010010011110011100011100" when "1000101110",
   "10001011110000000100110001001000000110001000100100001000111" when "1000101111",
   "10001100000000000100110010001110000001111101010101110100000" when "1000110000",
   "10001100010000000100110011010100000101110010001000100101001" when "1000110001",
   "10001100100000000100110100011010010001100110111100011100011" when "1000110010",
   "10001100110000000100110101100000100101011011110001011010000" when "1000110011",
   "10001101000000000100110110100111000001010000100111011101111" when "1000110100",
   "10001101010000000100110111101101100101000101011110101000010" when "1000110101",
   "10001101100000000100111000110100010000111010010110111001010" when "1000110110",
   "10001101110000000100111001111011000100101111010000010001000" when "1000110111",
   "10001110000000000100111011000010000000100100001010101111110" when "1000111000",
   "10001110010000000100111100001001000100011001000110010101011" when "1000111001",
   "10001110100000000100111101010000010000001110000011000010001" when "1000111010",
   "10001110110000000100111110010111100100000011000000110110001" when "1000111011",
   "10001111000000000100111111011110111111110111111111110001100" when "1000111100",
   "10001111010000000101000000100110100011101100111111110100011" when "1000111101",
   "10001111100000000101000001101110001111100010000000111110111" when "1000111110",
   "10001111110000000101000010110110000011010111000011010001001" when "1000111111",
   "10010000000000000101000011111101111111001100000110101011010" when "1001000000",
   "10010000010000000101000101000110000011000001001011001101011" when "1001000001",
   "10010000100000000101000110001110001110110110010000110111101" when "1001000010",
   "10010000110000000101000111010110100010101011010111101010001" when "1001000011",
   "10010001000000000101001000011110111110100000011111100101000" when "1001000100",
   "10010001010000000101001001100111100010010101101000101000011" when "1001000101",
   "10010001100000000101001010110000001110001010110010110100011" when "1001000110",
   "10010001110000000101001011111001000001111111111110001001001" when "1001000111",
   "10010010000000000101001101000001111101110101001010100110110" when "1001001000",
   "10010010010000000101001110001011000001101010011000001101011" when "1001001001",
   "10010010100000000101001111010100001101011111100110111101001" when "1001001010",
   "10010010110000000101010000011101100001010100110110110110000" when "1001001011",
   "10010011000000000101010001100110111101001010000111111000011" when "1001001100",
   "10010011010000000101010010110000100000111111011010000100010" when "1001001101",
   "10010011100000000101010011111010001100110100101101011001110" when "1001001110",
   "10010011110000000101010101000100000000101010000001111001000" when "1001001111",
   "10010100000000000101010110001101111100011111010111100010000" when "1001010000",
   "10010100010000000101010111011000000000010100101110010101001" when "1001010001",
   "10010100100000000101011000100010001100001010000110010010011" when "1001010010",
   "10010100110000000101011001101100011111111111011111011001111" when "1001010011",
   "10010101000000000101011010110110111011110100111001101011101" when "1001010100",
   "10010101010000000101011100000001011111101010010101001000000" when "1001010101",
   "10010101100000000101011101001100001011011111110001101111000" when "1001010110",
   "10010101110000000101011110010110111111010101001111100000101" when "1001010111",
   "10010110000000000101011111100001111011001010101110011101010" when "1001011000",
   "10010110010000000101100000101100111111000000001110100100111" when "1001011001",
   "10010110100000000101100001111000001010110101101111110111100" when "1001011010",
   "10010110110000000101100011000011011110101011010010010101100" when "1001011011",
   "10010111000000000101100100001110111010100000110101111110110" when "1001011100",
   "10010111010000000101100101011010011110010110011010110011101" when "1001011101",
   "10010111100000000101100110100110001010001100000000110100001" when "1001011110",
   "10010111110000000101100111110001111110000001101000000000010" when "1001011111",
   "10011000000000000101101000111101111001110111010000011000011" when "1001100000",
   "10011000010000000101101010001001111101101100111001111100011" when "1001100001",
   "10011000100000000101101011010110001001100010100100101100101" when "1001100010",
   "10011000110000000101101100100010011101011000010000101001000" when "1001100011",
   "10011001000000000101101101101110111001001101111101110001111" when "1001100100",
   "10011001010000000101101110111011011101000011101100000111001" when "1001100101",
   "10011001100000000101110000001000001000111001011011101001000" when "1001100110",
   "10011001110000000101110001010100111100101111001100010111110" when "1001100111",
   "10011010000000000101110010100001111000100100111110010011010" when "1001101000",
   "10011010010000000101110011101110111100011010110001011011111" when "1001101001",
   "10011010100000000101110100111100001000010000100101110001100" when "1001101010",
   "10011010110000000101110110001001011100000110011011010100011" when "1001101011",
   "10011011000000000101110111010110110111111100010010000100110" when "1001101100",
   "10011011010000000101111000100100011011110010001010000010100" when "1001101101",
   "10011011100000000101111001110010000111101000000011001101111" when "1001101110",
   "10011011110000000101111010111111111011011101111101100111001" when "1001101111",
   "10011100000000000101111100001101110111010011111001001110001" when "1001110000",
   "10011100010000000101111101011011111011001001110110000011001" when "1001110001",
   "10011100100000000101111110101010000110111111110100000110011" when "1001110010",
   "10011100110000000101111111111000011010110101110011010111110" when "1001110011",
   "10011101000000000110000001000110110110101011110011110111100" when "1001110100",
   "10011101010000000110000010010101011010100001110101100101110" when "1001110101",
   "10011101100000000110000011100100000110010111111000100010101" when "1001110110",
   "10011101110000000110000100110010111010001101111100101110011" when "1001110111",
   "10011110000000000110000110000001110110000100000010001000111" when "1001111000",
   "10011110010000000110000111010000111001111010001000110010011" when "1001111001",
   "10011110100000000110001000100000000101110000010000101011000" when "1001111010",
   "10011110110000000110001001101111011001100110011001110010111" when "1001111011",
   "10011111000000000110001010111110110101011100100100001010001" when "1001111100",
   "10011111010000000110001100001110011001010010101111110001000" when "1001111101",
   "10011111100000000110001101011110000101001000111100100111011" when "1001111110",
   "10011111110000000110001110101101111000111111001010101101100" when "1001111111",
   "10100000000000000110001111111101110100110101011010000011100" when "1010000000",
   "10100000010000000110010001001101111000101011101010101001100" when "1010000001",
   "10100000100000000110010010011110000100100001111100011111101" when "1010000010",
   "10100000110000000110010011101110011000011000001111100110000" when "1010000011",
   "10100001000000000110010100111110110100001110100011111100110" when "1010000100",
   "10100001010000000110010110001111011000000100111001100100000" when "1010000101",
   "10100001100000000110010111100000000011111011010000011011111" when "1010000110",
   "10100001110000000110011000110000110111110001101000100100100" when "1010000111",
   "10100010000000000110011010000001110011101000000001111110000" when "1010001000",
   "10100010010000000110011011010010110111011110011100101000100" when "1010001001",
   "10100010100000000110011100100100000011010100111000100100001" when "1010001010",
   "10100010110000000110011101110101010111001011010101110001000" when "1010001011",
   "10100011000000000110011111000110110011000001110100001111010" when "1010001100",
   "10100011010000000110100000011000010110111000010011111111000" when "1010001101",
   "10100011100000000110100001101010000010101110110101000000011" when "1010001110",
   "10100011110000000110100010111011110110100101010111010011100" when "1010001111",
   "10100100000000000110100100001101110010011011111010111000011" when "1010010000",
   "10100100010000000110100101011111110110010010011111101111011" when "1010010001",
   "10100100100000000110100110110010000010001001000101111000100" when "1010010010",
   "10100100110000000110101000000100010101111111101101010011111" when "1010010011",
   "10100101000000000110101001010110110001110110010110000001101" when "1010010100",
   "10100101010000000110101010101001010101101101000000000001111" when "1010010101",
   "10100101100000000110101011111100000001100011101011010100101" when "1010010110",
   "10100101110000000110101101001110110101011010010111111010010" when "1010010111",
   "10100110000000000110101110100001110001010001000101110010110" when "1010011000",
   "10100110010000000110101111110100110101000111110100111110010" when "1010011001",
   "10100110100000000110110001001000000000111110100101011100111" when "1010011010",
   "10100110110000000110110010011011010100110101010111001110101" when "1010011011",
   "10100111000000000110110011101110110000101100001010010011111" when "1010011100",
   "10100111010000000110110101000010010100100010111110101100101" when "1010011101",
   "10100111100000000110110110010110000000011001110100011000111" when "1010011110",
   "10100111110000000110110111101001110100010000101011011001000" when "1010011111",
   "10101000000000000110111000111101110000000111100011101101000" when "1010100000",
   "10101000010000000110111010010001110011111110011101010101000" when "1010100001",
   "10101000100000000110111011100101111111110101011000010001000" when "1010100010",
   "10101000110000000110111100111010010011101100010100100001011" when "1010100011",
   "10101001000000000110111110001110101111100011010010000110001" when "1010100100",
   "10101001010000000110111111100011010011011010010000111111010" when "1010100101",
   "10101001100000000111000000110111111111010001010001001101001" when "1010100110",
   "10101001110000000111000010001100110011001000010010101111101" when "1010100111",
   "10101010000000000111000011100001101110111111010101100111001" when "1010101000",
   "10101010010000000111000100110110110010110110011001110011101" when "1010101001",
   "10101010100000000111000110001011111110101101011111010101001" when "1010101010",
   "10101010110000000111000111100001010010100100100110001100000" when "1010101011",
   "10101011000000000111001000110110101110011011101110011000001" when "1010101100",
   "10101011010000000111001010001100010010010010110111111001111" when "1010101101",
   "10101011100000000111001011100001111110001010000010110001001" when "1010101110",
   "10101011110000000111001100110111110010000001001110111110010" when "1010101111",
   "10101100000000000111001110001101101101111000011100100001010" when "1010110000",
   "10101100010000000111001111100011110001101111101011011010001" when "1010110001",
   "10101100100000000111010000111001111101100110111011101001010" when "1010110010",
   "10101100110000000111010010010000010001011110001101001110100" when "1010110011",
   "10101101000000000111010011100110101101010101100000001010010" when "1010110100",
   "10101101010000000111010100111101010001001100110100011100011" when "1010110101",
   "10101101100000000111010110010011111101000100001010000101001" when "1010110110",
   "10101101110000000111010111101010110000111011100001000100110" when "1010110111",
   "10101110000000000111011001000001101100110010111001011011001" when "1010111000",
   "10101110010000000111011010011000110000101010010011001000101" when "1010111001",
   "10101110100000000111011011101111111100100001101110001101001" when "1010111010",
   "10101110110000000111011101000111010000011001001010101001000" when "1010111011",
   "10101111000000000111011110011110101100010000101000011100001" when "1010111100",
   "10101111010000000111011111110110010000001000000111100110110" when "1010111101",
   "10101111100000000111100001001101111011111111101000001001001" when "1010111110",
   "10101111110000000111100010100101101111110111001010000011001" when "1010111111",
   "10110000000000000111100011111101101011101110101101010101001" when "1011000000",
   "10110000010000000111100101010101101111100110010001111111000" when "1011000001",
   "10110000100000000111100110101101111011011101111000000001000" when "1011000010",
   "10110000110000000111101000000110001111010101011111011011011" when "1011000011",
   "10110001000000000111101001011110101011001101001000001110000" when "1011000100",
   "10110001010000000111101010110111001111000100110010011001001" when "1011000101",
   "10110001100000000111101100001111111010111100011101111101000" when "1011000110",
   "10110001110000000111101101101000101110110100001010111001100" when "1011000111",
   "10110010000000000111101111000001101010101011111001001110111" when "1011001000",
   "10110010010000000111110000011010101110100011101000111101011" when "1011001001",
   "10110010100000000111110001110011111010011011011010000100111" when "1011001010",
   "10110010110000000111110011001101001110010011001100100101101" when "1011001011",
   "10110011000000000111110100100110101010001011000000011111110" when "1011001100",
   "10110011010000000111110110000000001110000010110101110011100" when "1011001101",
   "10110011100000000111110111011001111001111010101100100000110" when "1011001110",
   "10110011110000000111111000110011101101110010100100100111110" when "1011001111",
   "10110100000000000111111010001101101001101010011110001000101" when "1011010000",
   "10110100010000000111111011100111101101100010011001000011101" when "1011010001",
   "10110100100000000111111101000001111001011010010101011000101" when "1011010010",
   "10110100110000000111111110011100001101010010010011000111111" when "1011010011",
   "10110101000000000111111111110110101001001010010010010001100" when "1011010100",
   "10110101010000001000000001010001001101000010010010110101101" when "1011010101",
   "10110101100000001000000010101011111000111010010100110100100" when "1011010110",
   "10110101110000001000000100000110101100110010011000001110000" when "1011010111",
   "10110110000000001000000101100001101000101010011101000010011" when "1011011000",
   "10110110010000001000000110111100101100100010100011010001110" when "1011011001",
   "10110110100000001000001000010111111000011010101010111100010" when "1011011010",
   "10110110110000001000001001110011001100010010110100000010000" when "1011011011",
   "10110111000000001000001011001110101000001010111110100011010" when "1011011100",
   "10110111010000001000001100101010001100000011001010011111111" when "1011011101",
   "10110111100000001000001110000101110111111011010111111000001" when "1011011110",
   "10110111110000001000001111100001101011110011100110101100001" when "1011011111",
   "10111000000000001000010000111101100111101011110110111100000" when "1011100000",
   "10111000010000001000010010011001101011100100001000100111111" when "1011100001",
   "10111000100000001000010011110101110111011100011011101111111" when "1011100010",
   "10111000110000001000010101010010001011010100110000010100001" when "1011100011",
   "10111001000000001000010110101110100111001101000110010100110" when "1011100100",
   "10111001010000001000011000001011001011000101011101110001111" when "1011100101",
   "10111001100000001000011001100111110110111101110110101011110" when "1011100110",
   "10111001110000001000011011000100101010110110010001000010010" when "1011100111",
   "10111010000000001000011100100001100110101110101100110101101" when "1011101000",
   "10111010010000001000011101111110101010100111001010000110000" when "1011101001",
   "10111010100000001000011111011011110110011111101000110011100" when "1011101010",
   "10111010110000001000100000111001001010011000001000111110010" when "1011101011",
   "10111011000000001000100010010110100110010000101010100110011" when "1011101100",
   "10111011010000001000100011110100001010001001001101101100000" when "1011101101",
   "10111011100000001000100101010001110110000001110010001111010" when "1011101110",
   "10111011110000001000100110101111101001111010011000010000010" when "1011101111",
   "10111100000000001000101000001101100101110010111111101111001" when "1011110000",
   "10111100010000001000101001101011101001101011101000101100000" when "1011110001",
   "10111100100000001000101011001001110101100100010011000111000" when "1011110010",
   "10111100110000001000101100101000001001011100111111000000010" when "1011110011",
   "10111101000000001000101110000110100101010101101100010111111" when "1011110100",
   "10111101010000001000101111100101001001001110011011001110000" when "1011110101",
   "10111101100000001000110001000011110101000111001011100010110" when "1011110110",
   "10111101110000001000110010100010101000111111111101010110010" when "1011110111",
   "10111110000000001000110100000001100100111000110000101000101" when "1011111000",
   "10111110010000001000110101100000101000110001100101011010000" when "1011111001",
   "10111110100000001000110110111111110100101010011011101010100" when "1011111010",
   "10111110110000001000111000011111001000100011010011011010010" when "1011111011",
   "10111111000000001000111001111110100100011100001100101001010" when "1011111100",
   "10111111010000001000111011011110001000010101000111010111111" when "1011111101",
   "10111111100000001000111100111101110100001110000011100110001" when "1011111110",
   "10111111110000001000111110011101101000000111000001010100001" when "1011111111",
   "11000000000000001000111111111101100100000000000000100010000" when "1100000000",
   "11000000010000001001000001011101100111111001000001001111111" when "1100000001",
   "11000000100000001001000010111101110011110010000011011101111" when "1100000010",
   "11000000110000001001000100011110000111101011000111001100001" when "1100000011",
   "11000001000000001001000101111110100011100100001100011010110" when "1100000100",
   "11000001010000001001000111011111000111011101010011001001111" when "1100000101",
   "11000001100000001001001000111111110011010110011011011001101" when "1100000110",
   "11000001110000001001001010100000100111001111100101001010000" when "1100000111",
   "11000010000000001001001100000001100011001000110000011011011" when "1100001000",
   "11000010010000001001001101100010100111000001111101001101110" when "1100001001",
   "11000010100000001001001111000011110010111011001011100001010" when "1100001010",
   "11000010110000001001010000100101000110110100011011010110000" when "1100001011",
   "11000011000000001001010010000110100010101101101100101100001" when "1100001100",
   "11000011010000001001010011101000000110100110111111100011110" when "1100001101",
   "11000011100000001001010101001001110010100000010011111101000" when "1100001110",
   "11000011110000001001010110101011100110011001101001110111111" when "1100001111",
   "11000100000000001001011000001101100010010011000001010100110" when "1100010000",
   "11000100010000001001011001101111100110001100011010010011101" when "1100010001",
   "11000100100000001001011011010001110010000101110100110100101" when "1100010010",
   "11000100110000001001011100110100000101111111010000110111111" when "1100010011",
   "11000101000000001001011110010110100001111000101110011101100" when "1100010100",
   "11000101010000001001011111111001000101110010001101100101100" when "1100010101",
   "11000101100000001001100001011011110001101011101110010000010" when "1100010110",
   "11000101110000001001100010111110100101100101010000011101110" when "1100010111",
   "11000110000000001001100100100001100001011110110100001110001" when "1100011000",
   "11000110010000001001100110000100100101011000011001100001100" when "1100011001",
   "11000110100000001001100111100111110001010010000000011000000" when "1100011010",
   "11000110110000001001101001001011000101001011101000110001101" when "1100011011",
   "11000111000000001001101010101110100001000101010010101110110" when "1100011100",
   "11000111010000001001101100010010000100111110111110001111011" when "1100011101",
   "11000111100000001001101101110101110000111000101011010011101" when "1100011110",
   "11000111110000001001101111011001100100110010011001111011101" when "1100011111",
   "11001000000000001001110000111101100000101100001010000111011" when "1100100000",
   "11001000010000001001110010100001100100100101111011110111010" when "1100100001",
   "11001000100000001001110100000101110000011111101111001011010" when "1100100010",
   "11001000110000001001110101101010000100011001100100000011100" when "1100100011",
   "11001001000000001001110111001110100000010011011010100000001" when "1100100100",
   "11001001010000001001111000110011000100001101010010100001001" when "1100100101",
   "11001001100000001001111010010111110000000111001100000110111" when "1100100110",
   "11001001110000001001111011111100100100000001000111010001011" when "1100100111",
   "11001010000000001001111101100001011111111011000100000000110" when "1100101000",
   "11001010010000001001111111000110100011110101000010010101000" when "1100101001",
   "11001010100000001010000000101011101111101111000010001110100" when "1100101010",
   "11001010110000001010000010010001000011101001000011101101010" when "1100101011",
   "11001011000000001010000011110110011111100011000110110001011" when "1100101100",
   "11001011010000001010000101011100000011011101001011011011000" when "1100101101",
   "11001011100000001010000111000001101111010111010001101010001" when "1100101110",
   "11001011110000001010001000100111100011010001011001011111001" when "1100101111",
   "11001100000000001010001010001101011111001011100010111010000" when "1100110000",
   "11001100010000001010001011110011100011000101101101111010111" when "1100110001",
   "11001100100000001010001101011001101110111111111010100001110" when "1100110010",
   "11001100110000001010001111000000000010111010001000101111000" when "1100110011",
   "11001101000000001010010000100110011110110100011000100010101" when "1100110100",
   "11001101010000001010010010001101000010101110101001111100110" when "1100110101",
   "11001101100000001010010011110011101110101000111100111101011" when "1100110110",
   "11001101110000001010010101011010100010100011010001100100111" when "1100110111",
   "11001110000000001010010111000001011110011101100111110011010" when "1100111000",
   "11001110010000001010011000101000100010010111111111101000101" when "1100111001",
   "11001110100000001010011010001111101110010010011001000101000" when "1100111010",
   "11001110110000001010011011110111000010001100110100001000110" when "1100111011",
   "11001111000000001010011101011110011110000111010000110011111" when "1100111100",
   "11001111010000001010011111000110000010000001101111000110100" when "1100111101",
   "11001111100000001010100000101101101101111100001111000000101" when "1100111110",
   "11001111110000001010100010010101100001110110110000100010101" when "1100111111",
   "11010000000000001010100011111101011101110001010011101100100" when "1101000000",
   "11010000010000001010100101100101100001101011111000011110011" when "1101000001",
   "11010000100000001010100111001101101101100110011110111000010" when "1101000010",
   "11010000110000001010101000110110000001100001000110111010100" when "1101000011",
   "11010001000000001010101010011110011101011011110000100101001" when "1101000100",
   "11010001010000001010101100000111000001010110011011111000010" when "1101000101",
   "11010001100000001010101101101111101101010001001000110011111" when "1101000110",
   "11010001110000001010101111011000100001001011110111011000011" when "1101000111",
   "11010010000000001010110001000001011101000110100111100101110" when "1101001000",
   "11010010010000001010110010101010100001000001011001011100001" when "1101001001",
   "11010010100000001010110100010011101100111100001100111011100" when "1101001010",
   "11010010110000001010110101111101000000110111000010000100010" when "1101001011",
   "11010011000000001010110111100110011100110001111000110110011" when "1101001100",
   "11010011010000001010111001010000000000101100110001010010000" when "1101001101",
   "11010011100000001010111010111001101100100111101011010111001" when "1101001110",
   "11010011110000001010111100100011100000100010100111000110001" when "1101001111",
   "11010100000000001010111110001101011100011101100100011111000" when "1101010000",
   "11010100010000001010111111110111100000011000100011100001111" when "1101010001",
   "11010100100000001011000001100001101100010011100100001110110" when "1101010010",
   "11010100110000001011000011001100000000001110100110100110000" when "1101010011",
   "11010101000000001011000100110110011100001001101010100111101" when "1101010100",
   "11010101010000001011000110100001000000000100110000010011110" when "1101010101",
   "11010101100000001011001000001011101011111111110111101010011" when "1101010110",
   "11010101110000001011001001110110011111111011000000101011111" when "1101010111",
   "11010110000000001011001011100001011011110110001011011000010" when "1101011000",
   "11010110010000001011001101001100011111110001010111101111101" when "1101011001",
   "11010110100000001011001110110111101011101100100101110010000" when "1101011010",
   "11010110110000001011010000100010111111100111110101011111110" when "1101011011",
   "11010111000000001011010010001110011011100011000110111000111" when "1101011100",
   "11010111010000001011010011111001111111011110011001111101100" when "1101011101",
   "11010111100000001011010101100101101011011001101110101101110" when "1101011110",
   "11010111110000001011010111010001011111010101000101001001101" when "1101011111",
   "11011000000000001011011000111101011011010000011101010001100" when "1101100000",
   "11011000010000001011011010101001011111001011110111000101011" when "1101100001",
   "11011000100000001011011100010101101011000111010010100101011" when "1101100010",
   "11011000110000001011011110000001111111000010101111110001100" when "1101100011",
   "11011001000000001011011111101110011010111110001110101010001" when "1101100100",
   "11011001010000001011100001011010111110111001101111001111010" when "1101100101",
   "11011001100000001011100011000111101010110101010001100001000" when "1101100110",
   "11011001110000001011100100110100011110110000110101011111100" when "1101100111",
   "11011010000000001011100110100001011010101100011011001010110" when "1101101000",
   "11011010010000001011101000001110011110101000000010100011001" when "1101101001",
   "11011010100000001011101001111011101010100011101011101000101" when "1101101010",
   "11011010110000001011101011101000111110011111010110011011011" when "1101101011",
   "11011011000000001011101101010110011010011011000010111011100" when "1101101100",
   "11011011010000001011101111000011111110010110110001001001000" when "1101101101",
   "11011011100000001011110000110001101010010010100001000100010" when "1101101110",
   "11011011110000001011110010011111011110001110010010101101010" when "1101101111",
   "11011100000000001011110100001101011010001010000110000100001" when "1101110000",
   "11011100010000001011110101111011011110000101111011001001000" when "1101110001",
   "11011100100000001011110111101001101010000001110001111100000" when "1101110010",
   "11011100110000001011111001010111111101111101101010011101001" when "1101110011",
   "11011101000000001011111011000110011001111001100100101100110" when "1101110100",
   "11011101010000001011111100110100111101110101100000101010111" when "1101110101",
   "11011101100000001011111110100011101001110001011110010111101" when "1101110110",
   "11011101110000001100000000010010011101101101011101110011001" when "1101110111",
   "11011110000000001100000010000001011001101001011110111101100" when "1101111000",
   "11011110010000001100000011110000011101100101100001110110110" when "1101111001",
   "11011110100000001100000101011111101001100001100110011111010" when "1101111010",
   "11011110110000001100000111001110111101011101101100110111000" when "1101111011",
   "11011111000000001100001000111110011001011001110100111110001" when "1101111100",
   "11011111010000001100001010101101111101010101111110110100110" when "1101111101",
   "11011111100000001100001100011101101001010010001010011011000" when "1101111110",
   "11011111110000001100001110001101011101001110010111110001000" when "1101111111",
   "11100000000000001100001111111101011001001010100110110110110" when "1110000000",
   "11100000010000001100010001101101011101000110110111101100101" when "1110000001",
   "11100000100000001100010011011101101001000011001010010010101" when "1110000010",
   "11100000110000001100010101001101111100111111011110101000111" when "1110000011",
   "11100001000000001100010110111110011000111011110100101111100" when "1110000100",
   "11100001010000001100011000101110111100111000001100100110101" when "1110000101",
   "11100001100000001100011010011111101000110100100110001110011" when "1110000110",
   "11100001110000001100011100010000011100110001000001100110111" when "1110000111",
   "11100010000000001100011110000001011000101101011110110000010" when "1110001000",
   "11100010010000001100011111110010011100101001111101101010101" when "1110001001",
   "11100010100000001100100001100011101000100110011110010110001" when "1110001010",
   "11100010110000001100100011010100111100100011000000110010111" when "1110001011",
   "11100011000000001100100101000110011000011111100101000000111" when "1110001100",
   "11100011010000001100100110110111111100011100001011000000100" when "1110001101",
   "11100011100000001100101000101001101000011000110010110001110" when "1110001110",
   "11100011110000001100101010011011011100010101011100010100110" when "1110001111",
   "11100100000000001100101100001101011000010010000111101001101" when "1110010000",
   "11100100010000001100101101111111011100001110110100110000100" when "1110010001",
   "11100100100000001100101111110001101000001011100011101001100" when "1110010010",
   "11100100110000001100110001100011111100001000010100010100110" when "1110010011",
   "11100101000000001100110011010110011000000101000110110010011" when "1110010100",
   "11100101010000001100110101001000111100000001111011000010100" when "1110010101",
   "11100101100000001100110110111011100111111110110001000101010" when "1110010110",
   "11100101110000001100111000101110011011111011101000111010110" when "1110010111",
   "11100110000000001100111010100001010111111000100010100011001" when "1110011000",
   "11100110010000001100111100010100011011110101011101111110100" when "1110011001",
   "11100110100000001100111110000111100111110010011011001101000" when "1110011010",
   "11100110110000001100111111111010111011101111011010001110110" when "1110011011",
   "11100111000000001101000001101110010111101100011011000011111" when "1110011100",
   "11100111010000001101000011100001111011101001011101101100100" when "1110011101",
   "11100111100000001101000101010101100111100110100010001000110" when "1110011110",
   "11100111110000001101000111001001011011100011101000011000111" when "1110011111",
   "11101000000000001101001000111101010111100000110000011100110" when "1110100000",
   "11101000010000001101001010110001011011011101111010010100101" when "1110100001",
   "11101000100000001101001100100101100111011011000110000000101" when "1110100010",
   "11101000110000001101001110011001111011011000010011100000111" when "1110100011",
   "11101001000000001101010000001110010111010101100010110101100" when "1110100100",
   "11101001010000001101010010000010111011010010110011111110101" when "1110100101",
   "11101001100000001101010011110111100111010000000110111100011" when "1110100110",
   "11101001110000001101010101101100011011001101011011101110111" when "1110100111",
   "11101010000000001101010111100001010111001010110010010110010" when "1110101000",
   "11101010010000001101011001010110011011001000001010110010110" when "1110101001",
   "11101010100000001101011011001011100111000101100101000100010" when "1110101010",
   "11101010110000001101011101000000111011000011000001001011000" when "1110101011",
   "11101011000000001101011110110110010111000000011111000111001" when "1110101100",
   "11101011010000001101100000101011111010111101111110111000110" when "1110101101",
   "11101011100000001101100010100001100110111011100000100000000" when "1110101110",
   "11101011110000001101100100010111011010111001000011111101001" when "1110101111",
   "11101100000000001101100110001101010110110110101001010000000" when "1110110000",
   "11101100010000001101101000000011011010110100010000011000111" when "1110110001",
   "11101100100000001101101001111001100110110001111001010111111" when "1110110010",
   "11101100110000001101101011101111111010101111100100001101001" when "1110110011",
   "11101101000000001101101101100110010110101101010000111000111" when "1110110100",
   "11101101010000001101101111011100111010101010111111011011000" when "1110110101",
   "11101101100000001101110001010011100110101000101111110011110" when "1110110110",
   "11101101110000001101110011001010011010100110100010000011010" when "1110110111",
   "11101110000000001101110101000001010110100100010110001001110" when "1110111000",
   "11101110010000001101110110111000011010100010001100000111001" when "1110111001",
   "11101110100000001101111000101111100110100000000011111011101" when "1110111010",
   "11101110110000001101111010100110111010011101111101100111100" when "1110111011",
   "11101111000000001101111100011110010110011011111001001010101" when "1110111100",
   "11101111010000001101111110010101111010011001110110100101010" when "1110111101",
   "11101111100000001110000000001101100110010111110101110111101" when "1110111110",
   "11101111110000001110000010000101011010010101110111000001101" when "1110111111",
   "11110000000000001110000011111101010110010011111010000011100" when "1111000000",
   "11110000010000001110000101110101011010010001111110111101100" when "1111000001",
   "11110000100000001110000111101101100110010000000101101111100" when "1111000010",
   "11110000110000001110001001100101111010001110001110011001110" when "1111000011",
   "11110001000000001110001011011110010110001100011000111100100" when "1111000100",
   "11110001010000001110001101010110111010001010100101010111101" when "1111000101",
   "11110001100000001110001111001111100110001000110011101011011" when "1111000110",
   "11110001110000001110010001001000011010000111000011111000000" when "1111000111",
   "11110010000000001110010011000001010110000101010101111101011" when "1111001000",
   "11110010010000001110010100111010011010000011101001111011111" when "1111001001",
   "11110010100000001110010110110011100110000001111111110011011" when "1111001010",
   "11110010110000001110011000101100111010000000010111100100010" when "1111001011",
   "11110011000000001110011010100110010101111110110001001110011" when "1111001100",
   "11110011010000001110011100011111111001111101001100110010001" when "1111001101",
   "11110011100000001110011110011001100101111011101010001111011" when "1111001110",
   "11110011110000001110100000010011011001111010001001100110100" when "1111001111",
   "11110100000000001110100010001101010101111000101010110111011" when "1111010000",
   "11110100010000001110100100000111011001110111001110000010011" when "1111010001",
   "11110100100000001110100110000001100101110101110011000111011" when "1111010010",
   "11110100110000001110100111111011111001110100011010000110110" when "1111010011",
   "11110101000000001110101001110110010101110011000011000000011" when "1111010100",
   "11110101010000001110101011110000111001110001101101110100101" when "1111010101",
   "11110101100000001110101101101011100101110000011010100011011" when "1111010110",
   "11110101110000001110101111100110011001101111001001001101000" when "1111010111",
   "11110110000000001110110001100001010101101101111001110001100" when "1111011000",
   "11110110010000001110110011011100011001101100101100010000111" when "1111011001",
   "11110110100000001110110101010111100101101011100000101011100" when "1111011010",
   "11110110110000001110110111010010111001101010010111000001011" when "1111011011",
   "11110111000000001110111001001110010101101001001111010010100" when "1111011100",
   "11110111010000001110111011001001111001101000001001011111010" when "1111011101",
   "11110111100000001110111101000101100101100111000101100111101" when "1111011110",
   "11110111110000001110111111000001011001100110000011101011101" when "1111011111",
   "11111000000000001111000000111101010101100101000011101011101" when "1111100000",
   "11111000010000001111000010111001011001100100000101100111101" when "1111100001",
   "11111000100000001111000100110101100101100011001001011111101" when "1111100010",
   "11111000110000001111000110110001111001100010001111010100000" when "1111100011",
   "11111001000000001111001000101110010101100001010111000100110" when "1111100100",
   "11111001010000001111001010101010111001100000100000110010000" when "1111100101",
   "11111001100000001111001100100111100101011111101100011011110" when "1111100110",
   "11111001110000001111001110100100011001011110111010000010011" when "1111100111",
   "11111010000000001111010000100001010101011110001001100101111" when "1111101000",
   "11111010010000001111010010011110011001011101011011000110011" when "1111101001",
   "11111010100000001111010100011011100101011100101110100100000" when "1111101010",
   "11111010110000001111010110011000111001011100000011111110111" when "1111101011",
   "11111011000000001111011000010110010101011011011011010111000" when "1111101100",
   "11111011010000001111011010010011111001011010110100101100110" when "1111101101",
   "11111011100000001111011100010001100101011010010000000000001" when "1111101110",
   "11111011110000001111011110001111011001011001101101010001010" when "1111101111",
   "11111100000000001111100000001101010101011001001100100000010" when "1111110000",
   "11111100010000001111100010001011011001011000101101101101010" when "1111110001",
   "11111100100000001111100100001001100101011000010000111000011" when "1111110010",
   "11111100110000001111100110000111111001010111110110000001110" when "1111110011",
   "11111101000000001111101000000110010101010111011101001001100" when "1111110100",
   "11111101010000001111101010000100111001010111000110001111110" when "1111110101",
   "11111101100000001111101100000011100101010110110001010100101" when "1111110110",
   "11111101110000001111101110000010011001010110011110011000010" when "1111110111",
   "11111110000000001111110000000001010101010110001101011010110" when "1111111000",
   "11111110010000001111110010000000011001010101111110011100010" when "1111111001",
   "11111110100000001111110011111111100101010101110001011100111" when "1111111010",
   "11111110110000001111110101111110111001010101100110011100110" when "1111111011",
   "11111111000000001111110111111110010101010101011101011100000" when "1111111100",
   "11111111010000001111111001111101111001010101010110011010110" when "1111111101",
   "11111111100000001111111011111101100101010101010001011001001" when "1111111110",
   "11111111110000001111111101111101011001010101001110010111011" when "1111111111",
   "-----------------------------------------------------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_74_f400_uid92
--                    (IntAdderAlternative_74_F400_uid96)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_74_f400_uid92 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(73 downto 0);
          Y : in  std_logic_vector(73 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(73 downto 0)   );
end entity;

architecture arch of IntAdder_74_f400_uid92 is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(32 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(31 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(32 downto 0);
signal sum_l1_idx1 :  std_logic_vector(31 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(73 downto 42)) + ( "0" & Y(73 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
   sum_l0_idx1 <= s_sum_l0_idx1(31 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(32 downto 32);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(31 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(32 downto 32);
   R <= sum_l1_idx1(31 downto 0) & sum_l0_idx0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_74_f400_uid100
--                    (IntAdderAlternative_74_F400_uid104)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_74_f400_uid100 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(73 downto 0);
          Y : in  std_logic_vector(73 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(73 downto 0)   );
end entity;

architecture arch of IntAdder_74_f400_uid100 is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(32 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(31 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(32 downto 0);
signal sum_l1_idx1 :  std_logic_vector(31 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(73 downto 42)) + ( "0" & Y(73 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
   sum_l0_idx1 <= s_sum_l0_idx1(31 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(32 downto 32);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(31 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(32 downto 32);
   R <= sum_l1_idx1(31 downto 0) & sum_l0_idx0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--              KCMTable_6_780414346020670_unsigned_F400_uid110
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity KCMTable_6_780414346020670_unsigned_F400_uid110 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of KCMTable_6_780414346020670_unsigned_F400_uid110 is
signal TableOut :  std_logic_vector(55 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "00000000000000000000000000000000000000000000000000000000" when "000000",
   "00000010110001011100100001011111110111110100011100111110" when "000001",
   "00000101100010111001000010111111101111101000111001111100" when "000010",
   "00001000010100010101100100011111100111011101010110111010" when "000011",
   "00001011000101110010000101111111011111010001110011111000" when "000100",
   "00001101110111001110100111011111010111000110010000110110" when "000101",
   "00010000101000101011001000111111001110111010101101110100" when "000110",
   "00010011011010000111101010011111000110101111001010110010" when "000111",
   "00010110001011100100001011111110111110100011100111110000" when "001000",
   "00011000111101000000101101011110110110011000000100101110" when "001001",
   "00011011101110011101001110111110101110001100100001101100" when "001010",
   "00011110011111111001110000011110100110000000111110101010" when "001011",
   "00100001010001010110010001111110011101110101011011101000" when "001100",
   "00100100000010110010110011011110010101101001111000100110" when "001101",
   "00100110110100001111010100111110001101011110010101100100" when "001110",
   "00101001100101101011110110011110000101010010110010100010" when "001111",
   "00101100010111001000010111111101111101000111001111100000" when "010000",
   "00101111001000100100111001011101110100111011101100011110" when "010001",
   "00110001111010000001011010111101101100110000001001011100" when "010010",
   "00110100101011011101111100011101100100100100100110011010" when "010011",
   "00110111011100111010011101111101011100011001000011011000" when "010100",
   "00111010001110010110111111011101010100001101100000010110" when "010101",
   "00111100111111110011100000111101001100000001111101010100" when "010110",
   "00111111110001010000000010011101000011110110011010010010" when "010111",
   "01000010100010101100100011111100111011101010110111010000" when "011000",
   "01000101010100001001000101011100110011011111010100001110" when "011001",
   "01001000000101100101100110111100101011010011110001001100" when "011010",
   "01001010110111000010001000011100100011001000001110001010" when "011011",
   "01001101101000011110101001111100011010111100101011001000" when "011100",
   "01010000011001111011001011011100010010110001001000000110" when "011101",
   "01010011001011010111101100111100001010100101100101000100" when "011110",
   "01010101111100110100001110011100000010011010000010000010" when "011111",
   "01011000101110010000101111111011111010001110011111000000" when "100000",
   "01011011011111101101010001011011110010000010111011111110" when "100001",
   "01011110010001001001110010111011101001110111011000111100" when "100010",
   "01100001000010100110010100011011100001101011110101111010" when "100011",
   "01100011110100000010110101111011011001100000010010111000" when "100100",
   "01100110100101011111010111011011010001010100101111110110" when "100101",
   "01101001010110111011111000111011001001001001001100110100" when "100110",
   "01101100001000011000011010011011000000111101101001110010" when "100111",
   "01101110111001110100111011111010111000110010000110110000" when "101000",
   "01110001101011010001011101011010110000100110100011101110" when "101001",
   "01110100011100101101111110111010101000011011000000101100" when "101010",
   "01110111001110001010100000011010100000001111011101101010" when "101011",
   "01111001111111100111000001111010011000000011111010101000" when "101100",
   "01111100110001000011100011011010001111111000010111100110" when "101101",
   "01111111100010100000000100111010000111101100110100100100" when "101110",
   "10000010010011111100100110011001111111100001010001100010" when "101111",
   "10000101000101011001000111111001110111010101101110100000" when "110000",
   "10000111110110110101101001011001101111001010001011011110" when "110001",
   "10001010101000010010001010111001100110111110101000011100" when "110010",
   "10001101011001101110101100011001011110110011000101011010" when "110011",
   "10010000001011001011001101111001010110100111100010011000" when "110100",
   "10010010111100100111101111011001001110011011111111010110" when "110101",
   "10010101101110000100010000111001000110010000011100010100" when "110110",
   "10011000011111100000110010011000111110000100111001010010" when "110111",
   "10011011010000111101010011111000110101111001010110010000" when "111000",
   "10011110000010011001110101011000101101101101110011001110" when "111001",
   "10100000110011110110010110111000100101100010010000001100" when "111010",
   "10100011100101010010111000011000011101010110101101001010" when "111011",
   "10100110010110101111011001111000010101001011001010001000" when "111100",
   "10101001001000001011111011011000001100111111100111000110" when "111101",
   "10101011111001101000011100111000000100110100000100000100" when "111110",
   "10101110101011000100111110010111111100101000100001000010" when "111111",
   "--------------------------------------------------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--              KCMTable_4_780414346020670_unsigned_F400_uid112
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity KCMTable_4_780414346020670_unsigned_F400_uid112 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(3 downto 0);
          Y : out  std_logic_vector(53 downto 0)   );
end entity;

architecture arch of KCMTable_4_780414346020670_unsigned_F400_uid112 is
signal TableOut :  std_logic_vector(53 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "000000000000000000000000000000000000000000000000000000" when "0000",
   "000010110001011100100001011111110111110100011100111110" when "0001",
   "000101100010111001000010111111101111101000111001111100" when "0010",
   "001000010100010101100100011111100111011101010110111010" when "0011",
   "001011000101110010000101111111011111010001110011111000" when "0100",
   "001101110111001110100111011111010111000110010000110110" when "0101",
   "010000101000101011001000111111001110111010101101110100" when "0110",
   "010011011010000111101010011111000110101111001010110010" when "0111",
   "010110001011100100001011111110111110100011100111110000" when "1000",
   "011000111101000000101101011110110110011000000100101110" when "1001",
   "011011101110011101001110111110101110001100100001101100" when "1010",
   "011110011111111001110000011110100110000000111110101010" when "1011",
   "100001010001010110010001111110011101110101011011101000" when "1100",
   "100100000010110010110011011110010101101001111000100110" when "1101",
   "100110110100001111010100111110001101011110010101100100" when "1110",
   "101001100101101011110110011110000101010010110010100010" when "1111",
   "------------------------------------------------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_61_f400_uid178
--                    (IntAdderAlternative_61_F400_uid182)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_61_f400_uid178 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(60 downto 0);
          Y : in  std_logic_vector(60 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(60 downto 0)   );
end entity;

architecture arch of IntAdder_61_f400_uid178 is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(19 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(18 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(19 downto 0);
signal sum_l1_idx1 :  std_logic_vector(18 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(60 downto 42)) + ( "0" & Y(60 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
   sum_l0_idx1 <= s_sum_l0_idx1(18 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(19 downto 19);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(18 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(19 downto 19);
   R <= sum_l1_idx1(18 downto 0) & sum_l0_idx0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--             IntIntKCM_16_780414346020670_unsigned_F400_uid108
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2009,2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntIntKCM_16_780414346020670_unsigned_F400_uid108 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(15 downto 0);
          R : out  std_logic_vector(65 downto 0)   );
end entity;

architecture arch of IntIntKCM_16_780414346020670_unsigned_F400_uid108 is
   component KCMTable_6_780414346020670_unsigned_F400_uid110 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(55 downto 0)   );
   end component;

   component KCMTable_4_780414346020670_unsigned_F400_uid112 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(3 downto 0);
             Y : out  std_logic_vector(53 downto 0)   );
   end component;

   component IntAdder_61_f400_uid178 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(60 downto 0);
             Y : in  std_logic_vector(60 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(60 downto 0)   );
   end component;

   component Compressor_23_3 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             X1 : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

signal d0 :  std_logic_vector(5 downto 0);
signal pp0 :  std_logic_vector(55 downto 0);
signal d1 :  std_logic_vector(5 downto 0);
signal pp1 :  std_logic_vector(55 downto 0);
signal d2 :  std_logic_vector(3 downto 0);
signal pp2 :  std_logic_vector(53 downto 0);
signal heap_bh119_w0_0 :  std_logic;
signal heap_bh119_w1_0 :  std_logic;
signal heap_bh119_w2_0 :  std_logic;
signal heap_bh119_w3_0 :  std_logic;
signal heap_bh119_w4_0 :  std_logic;
signal heap_bh119_w5_0 :  std_logic;
signal heap_bh119_w6_0, heap_bh119_w6_0_d1, heap_bh119_w6_0_d2 :  std_logic;
signal heap_bh119_w7_0, heap_bh119_w7_0_d1, heap_bh119_w7_0_d2 :  std_logic;
signal heap_bh119_w8_0, heap_bh119_w8_0_d1, heap_bh119_w8_0_d2 :  std_logic;
signal heap_bh119_w9_0, heap_bh119_w9_0_d1, heap_bh119_w9_0_d2 :  std_logic;
signal heap_bh119_w10_0, heap_bh119_w10_0_d1, heap_bh119_w10_0_d2 :  std_logic;
signal heap_bh119_w11_0, heap_bh119_w11_0_d1, heap_bh119_w11_0_d2 :  std_logic;
signal heap_bh119_w12_0 :  std_logic;
signal heap_bh119_w13_0, heap_bh119_w13_0_d1, heap_bh119_w13_0_d2 :  std_logic;
signal heap_bh119_w14_0 :  std_logic;
signal heap_bh119_w15_0, heap_bh119_w15_0_d1, heap_bh119_w15_0_d2 :  std_logic;
signal heap_bh119_w16_0 :  std_logic;
signal heap_bh119_w17_0, heap_bh119_w17_0_d1, heap_bh119_w17_0_d2 :  std_logic;
signal heap_bh119_w18_0 :  std_logic;
signal heap_bh119_w19_0, heap_bh119_w19_0_d1, heap_bh119_w19_0_d2 :  std_logic;
signal heap_bh119_w20_0 :  std_logic;
signal heap_bh119_w21_0, heap_bh119_w21_0_d1, heap_bh119_w21_0_d2 :  std_logic;
signal heap_bh119_w22_0 :  std_logic;
signal heap_bh119_w23_0, heap_bh119_w23_0_d1, heap_bh119_w23_0_d2 :  std_logic;
signal heap_bh119_w24_0 :  std_logic;
signal heap_bh119_w25_0, heap_bh119_w25_0_d1, heap_bh119_w25_0_d2 :  std_logic;
signal heap_bh119_w26_0 :  std_logic;
signal heap_bh119_w27_0, heap_bh119_w27_0_d1, heap_bh119_w27_0_d2 :  std_logic;
signal heap_bh119_w28_0 :  std_logic;
signal heap_bh119_w29_0, heap_bh119_w29_0_d1, heap_bh119_w29_0_d2 :  std_logic;
signal heap_bh119_w30_0 :  std_logic;
signal heap_bh119_w31_0, heap_bh119_w31_0_d1, heap_bh119_w31_0_d2 :  std_logic;
signal heap_bh119_w32_0 :  std_logic;
signal heap_bh119_w33_0, heap_bh119_w33_0_d1, heap_bh119_w33_0_d2 :  std_logic;
signal heap_bh119_w34_0 :  std_logic;
signal heap_bh119_w35_0, heap_bh119_w35_0_d1, heap_bh119_w35_0_d2 :  std_logic;
signal heap_bh119_w36_0 :  std_logic;
signal heap_bh119_w37_0, heap_bh119_w37_0_d1, heap_bh119_w37_0_d2 :  std_logic;
signal heap_bh119_w38_0 :  std_logic;
signal heap_bh119_w39_0, heap_bh119_w39_0_d1, heap_bh119_w39_0_d2 :  std_logic;
signal heap_bh119_w40_0 :  std_logic;
signal heap_bh119_w41_0, heap_bh119_w41_0_d1, heap_bh119_w41_0_d2 :  std_logic;
signal heap_bh119_w42_0 :  std_logic;
signal heap_bh119_w43_0, heap_bh119_w43_0_d1, heap_bh119_w43_0_d2 :  std_logic;
signal heap_bh119_w44_0 :  std_logic;
signal heap_bh119_w45_0, heap_bh119_w45_0_d1, heap_bh119_w45_0_d2 :  std_logic;
signal heap_bh119_w46_0 :  std_logic;
signal heap_bh119_w47_0, heap_bh119_w47_0_d1, heap_bh119_w47_0_d2 :  std_logic;
signal heap_bh119_w48_0 :  std_logic;
signal heap_bh119_w49_0, heap_bh119_w49_0_d1, heap_bh119_w49_0_d2 :  std_logic;
signal heap_bh119_w50_0 :  std_logic;
signal heap_bh119_w51_0, heap_bh119_w51_0_d1, heap_bh119_w51_0_d2 :  std_logic;
signal heap_bh119_w52_0 :  std_logic;
signal heap_bh119_w53_0, heap_bh119_w53_0_d1, heap_bh119_w53_0_d2 :  std_logic;
signal heap_bh119_w54_0 :  std_logic;
signal heap_bh119_w55_0, heap_bh119_w55_0_d1, heap_bh119_w55_0_d2 :  std_logic;
signal heap_bh119_w6_1, heap_bh119_w6_1_d1, heap_bh119_w6_1_d2 :  std_logic;
signal heap_bh119_w7_1, heap_bh119_w7_1_d1, heap_bh119_w7_1_d2 :  std_logic;
signal heap_bh119_w8_1, heap_bh119_w8_1_d1, heap_bh119_w8_1_d2 :  std_logic;
signal heap_bh119_w9_1, heap_bh119_w9_1_d1, heap_bh119_w9_1_d2 :  std_logic;
signal heap_bh119_w10_1, heap_bh119_w10_1_d1, heap_bh119_w10_1_d2 :  std_logic;
signal heap_bh119_w11_1, heap_bh119_w11_1_d1, heap_bh119_w11_1_d2 :  std_logic;
signal heap_bh119_w12_1 :  std_logic;
signal heap_bh119_w13_1 :  std_logic;
signal heap_bh119_w14_1 :  std_logic;
signal heap_bh119_w15_1 :  std_logic;
signal heap_bh119_w16_1 :  std_logic;
signal heap_bh119_w17_1 :  std_logic;
signal heap_bh119_w18_1 :  std_logic;
signal heap_bh119_w19_1 :  std_logic;
signal heap_bh119_w20_1 :  std_logic;
signal heap_bh119_w21_1 :  std_logic;
signal heap_bh119_w22_1 :  std_logic;
signal heap_bh119_w23_1 :  std_logic;
signal heap_bh119_w24_1 :  std_logic;
signal heap_bh119_w25_1 :  std_logic;
signal heap_bh119_w26_1 :  std_logic;
signal heap_bh119_w27_1 :  std_logic;
signal heap_bh119_w28_1 :  std_logic;
signal heap_bh119_w29_1 :  std_logic;
signal heap_bh119_w30_1 :  std_logic;
signal heap_bh119_w31_1 :  std_logic;
signal heap_bh119_w32_1 :  std_logic;
signal heap_bh119_w33_1 :  std_logic;
signal heap_bh119_w34_1 :  std_logic;
signal heap_bh119_w35_1 :  std_logic;
signal heap_bh119_w36_1 :  std_logic;
signal heap_bh119_w37_1 :  std_logic;
signal heap_bh119_w38_1 :  std_logic;
signal heap_bh119_w39_1 :  std_logic;
signal heap_bh119_w40_1 :  std_logic;
signal heap_bh119_w41_1 :  std_logic;
signal heap_bh119_w42_1 :  std_logic;
signal heap_bh119_w43_1 :  std_logic;
signal heap_bh119_w44_1 :  std_logic;
signal heap_bh119_w45_1 :  std_logic;
signal heap_bh119_w46_1 :  std_logic;
signal heap_bh119_w47_1 :  std_logic;
signal heap_bh119_w48_1 :  std_logic;
signal heap_bh119_w49_1 :  std_logic;
signal heap_bh119_w50_1 :  std_logic;
signal heap_bh119_w51_1 :  std_logic;
signal heap_bh119_w52_1 :  std_logic;
signal heap_bh119_w53_1 :  std_logic;
signal heap_bh119_w54_1 :  std_logic;
signal heap_bh119_w55_1 :  std_logic;
signal heap_bh119_w56_0 :  std_logic;
signal heap_bh119_w57_0 :  std_logic;
signal heap_bh119_w58_0, heap_bh119_w58_0_d1 :  std_logic;
signal heap_bh119_w59_0, heap_bh119_w59_0_d1 :  std_logic;
signal heap_bh119_w60_0, heap_bh119_w60_0_d1 :  std_logic;
signal heap_bh119_w61_0, heap_bh119_w61_0_d1 :  std_logic;
signal heap_bh119_w12_2 :  std_logic;
signal heap_bh119_w13_2 :  std_logic;
signal heap_bh119_w14_2 :  std_logic;
signal heap_bh119_w15_2 :  std_logic;
signal heap_bh119_w16_2 :  std_logic;
signal heap_bh119_w17_2 :  std_logic;
signal heap_bh119_w18_2 :  std_logic;
signal heap_bh119_w19_2 :  std_logic;
signal heap_bh119_w20_2 :  std_logic;
signal heap_bh119_w21_2 :  std_logic;
signal heap_bh119_w22_2 :  std_logic;
signal heap_bh119_w23_2 :  std_logic;
signal heap_bh119_w24_2 :  std_logic;
signal heap_bh119_w25_2 :  std_logic;
signal heap_bh119_w26_2 :  std_logic;
signal heap_bh119_w27_2 :  std_logic;
signal heap_bh119_w28_2 :  std_logic;
signal heap_bh119_w29_2 :  std_logic;
signal heap_bh119_w30_2 :  std_logic;
signal heap_bh119_w31_2 :  std_logic;
signal heap_bh119_w32_2 :  std_logic;
signal heap_bh119_w33_2 :  std_logic;
signal heap_bh119_w34_2 :  std_logic;
signal heap_bh119_w35_2 :  std_logic;
signal heap_bh119_w36_2 :  std_logic;
signal heap_bh119_w37_2 :  std_logic;
signal heap_bh119_w38_2 :  std_logic;
signal heap_bh119_w39_2 :  std_logic;
signal heap_bh119_w40_2 :  std_logic;
signal heap_bh119_w41_2 :  std_logic;
signal heap_bh119_w42_2 :  std_logic;
signal heap_bh119_w43_2 :  std_logic;
signal heap_bh119_w44_2 :  std_logic;
signal heap_bh119_w45_2 :  std_logic;
signal heap_bh119_w46_2 :  std_logic;
signal heap_bh119_w47_2 :  std_logic;
signal heap_bh119_w48_2 :  std_logic;
signal heap_bh119_w49_2 :  std_logic;
signal heap_bh119_w50_2 :  std_logic;
signal heap_bh119_w51_2 :  std_logic;
signal heap_bh119_w52_2 :  std_logic;
signal heap_bh119_w53_2 :  std_logic;
signal heap_bh119_w54_2 :  std_logic;
signal heap_bh119_w55_2 :  std_logic;
signal heap_bh119_w56_1 :  std_logic;
signal heap_bh119_w57_1 :  std_logic;
signal heap_bh119_w58_1, heap_bh119_w58_1_d1 :  std_logic;
signal heap_bh119_w59_1, heap_bh119_w59_1_d1 :  std_logic;
signal heap_bh119_w60_1, heap_bh119_w60_1_d1 :  std_logic;
signal heap_bh119_w61_1, heap_bh119_w61_1_d1 :  std_logic;
signal heap_bh119_w62_0, heap_bh119_w62_0_d1, heap_bh119_w62_0_d2 :  std_logic;
signal heap_bh119_w63_0, heap_bh119_w63_0_d1, heap_bh119_w63_0_d2 :  std_logic;
signal heap_bh119_w64_0, heap_bh119_w64_0_d1, heap_bh119_w64_0_d2 :  std_logic;
signal heap_bh119_w65_0, heap_bh119_w65_0_d1, heap_bh119_w65_0_d2 :  std_logic;
signal tempR_bh119_0, tempR_bh119_0_d1, tempR_bh119_0_d2, tempR_bh119_0_d3 :  std_logic_vector(5 downto 0);
signal CompressorIn_bh119_0_0 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_0_1 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_0_0 :  std_logic_vector(2 downto 0);
signal heap_bh119_w12_3, heap_bh119_w12_3_d1, heap_bh119_w12_3_d2 :  std_logic;
signal heap_bh119_w13_3, heap_bh119_w13_3_d1, heap_bh119_w13_3_d2 :  std_logic;
signal heap_bh119_w14_3, heap_bh119_w14_3_d1, heap_bh119_w14_3_d2 :  std_logic;
signal CompressorIn_bh119_1_2 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_1_3 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_1_1 :  std_logic_vector(2 downto 0);
signal heap_bh119_w14_4, heap_bh119_w14_4_d1, heap_bh119_w14_4_d2 :  std_logic;
signal heap_bh119_w15_3, heap_bh119_w15_3_d1, heap_bh119_w15_3_d2 :  std_logic;
signal heap_bh119_w16_3, heap_bh119_w16_3_d1, heap_bh119_w16_3_d2 :  std_logic;
signal CompressorIn_bh119_2_4 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_2_5 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_2_2 :  std_logic_vector(2 downto 0);
signal heap_bh119_w16_4, heap_bh119_w16_4_d1, heap_bh119_w16_4_d2 :  std_logic;
signal heap_bh119_w17_3, heap_bh119_w17_3_d1, heap_bh119_w17_3_d2 :  std_logic;
signal heap_bh119_w18_3, heap_bh119_w18_3_d1, heap_bh119_w18_3_d2 :  std_logic;
signal CompressorIn_bh119_3_6 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_3_7 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_3_3 :  std_logic_vector(2 downto 0);
signal heap_bh119_w18_4, heap_bh119_w18_4_d1, heap_bh119_w18_4_d2 :  std_logic;
signal heap_bh119_w19_3, heap_bh119_w19_3_d1, heap_bh119_w19_3_d2 :  std_logic;
signal heap_bh119_w20_3, heap_bh119_w20_3_d1, heap_bh119_w20_3_d2 :  std_logic;
signal CompressorIn_bh119_4_8 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_4_9 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_4_4 :  std_logic_vector(2 downto 0);
signal heap_bh119_w20_4, heap_bh119_w20_4_d1, heap_bh119_w20_4_d2 :  std_logic;
signal heap_bh119_w21_3, heap_bh119_w21_3_d1, heap_bh119_w21_3_d2 :  std_logic;
signal heap_bh119_w22_3, heap_bh119_w22_3_d1, heap_bh119_w22_3_d2 :  std_logic;
signal CompressorIn_bh119_5_10 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_5_11 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_5_5 :  std_logic_vector(2 downto 0);
signal heap_bh119_w22_4, heap_bh119_w22_4_d1, heap_bh119_w22_4_d2 :  std_logic;
signal heap_bh119_w23_3, heap_bh119_w23_3_d1, heap_bh119_w23_3_d2 :  std_logic;
signal heap_bh119_w24_3, heap_bh119_w24_3_d1, heap_bh119_w24_3_d2 :  std_logic;
signal CompressorIn_bh119_6_12 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_6_13 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_6_6 :  std_logic_vector(2 downto 0);
signal heap_bh119_w24_4, heap_bh119_w24_4_d1, heap_bh119_w24_4_d2 :  std_logic;
signal heap_bh119_w25_3, heap_bh119_w25_3_d1, heap_bh119_w25_3_d2 :  std_logic;
signal heap_bh119_w26_3, heap_bh119_w26_3_d1, heap_bh119_w26_3_d2 :  std_logic;
signal CompressorIn_bh119_7_14 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_7_15 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_7_7 :  std_logic_vector(2 downto 0);
signal heap_bh119_w26_4, heap_bh119_w26_4_d1, heap_bh119_w26_4_d2 :  std_logic;
signal heap_bh119_w27_3, heap_bh119_w27_3_d1, heap_bh119_w27_3_d2 :  std_logic;
signal heap_bh119_w28_3, heap_bh119_w28_3_d1, heap_bh119_w28_3_d2 :  std_logic;
signal CompressorIn_bh119_8_16 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_8_17 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_8_8 :  std_logic_vector(2 downto 0);
signal heap_bh119_w28_4, heap_bh119_w28_4_d1, heap_bh119_w28_4_d2 :  std_logic;
signal heap_bh119_w29_3, heap_bh119_w29_3_d1, heap_bh119_w29_3_d2 :  std_logic;
signal heap_bh119_w30_3, heap_bh119_w30_3_d1, heap_bh119_w30_3_d2 :  std_logic;
signal CompressorIn_bh119_9_18 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_9_19 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_9_9 :  std_logic_vector(2 downto 0);
signal heap_bh119_w30_4, heap_bh119_w30_4_d1, heap_bh119_w30_4_d2 :  std_logic;
signal heap_bh119_w31_3, heap_bh119_w31_3_d1, heap_bh119_w31_3_d2 :  std_logic;
signal heap_bh119_w32_3, heap_bh119_w32_3_d1, heap_bh119_w32_3_d2 :  std_logic;
signal CompressorIn_bh119_10_20 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_10_21 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_10_10 :  std_logic_vector(2 downto 0);
signal heap_bh119_w32_4, heap_bh119_w32_4_d1, heap_bh119_w32_4_d2 :  std_logic;
signal heap_bh119_w33_3, heap_bh119_w33_3_d1, heap_bh119_w33_3_d2 :  std_logic;
signal heap_bh119_w34_3, heap_bh119_w34_3_d1, heap_bh119_w34_3_d2 :  std_logic;
signal CompressorIn_bh119_11_22 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_11_23 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_11_11 :  std_logic_vector(2 downto 0);
signal heap_bh119_w34_4, heap_bh119_w34_4_d1, heap_bh119_w34_4_d2 :  std_logic;
signal heap_bh119_w35_3, heap_bh119_w35_3_d1, heap_bh119_w35_3_d2 :  std_logic;
signal heap_bh119_w36_3, heap_bh119_w36_3_d1, heap_bh119_w36_3_d2 :  std_logic;
signal CompressorIn_bh119_12_24 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_12_25 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_12_12 :  std_logic_vector(2 downto 0);
signal heap_bh119_w36_4, heap_bh119_w36_4_d1, heap_bh119_w36_4_d2 :  std_logic;
signal heap_bh119_w37_3, heap_bh119_w37_3_d1, heap_bh119_w37_3_d2 :  std_logic;
signal heap_bh119_w38_3, heap_bh119_w38_3_d1, heap_bh119_w38_3_d2 :  std_logic;
signal CompressorIn_bh119_13_26 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_13_27 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_13_13 :  std_logic_vector(2 downto 0);
signal heap_bh119_w38_4, heap_bh119_w38_4_d1, heap_bh119_w38_4_d2 :  std_logic;
signal heap_bh119_w39_3, heap_bh119_w39_3_d1, heap_bh119_w39_3_d2 :  std_logic;
signal heap_bh119_w40_3, heap_bh119_w40_3_d1, heap_bh119_w40_3_d2 :  std_logic;
signal CompressorIn_bh119_14_28 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_14_29 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_14_14 :  std_logic_vector(2 downto 0);
signal heap_bh119_w40_4, heap_bh119_w40_4_d1, heap_bh119_w40_4_d2 :  std_logic;
signal heap_bh119_w41_3, heap_bh119_w41_3_d1, heap_bh119_w41_3_d2 :  std_logic;
signal heap_bh119_w42_3, heap_bh119_w42_3_d1, heap_bh119_w42_3_d2 :  std_logic;
signal CompressorIn_bh119_15_30 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_15_31 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_15_15 :  std_logic_vector(2 downto 0);
signal heap_bh119_w42_4, heap_bh119_w42_4_d1, heap_bh119_w42_4_d2 :  std_logic;
signal heap_bh119_w43_3, heap_bh119_w43_3_d1, heap_bh119_w43_3_d2 :  std_logic;
signal heap_bh119_w44_3, heap_bh119_w44_3_d1, heap_bh119_w44_3_d2 :  std_logic;
signal CompressorIn_bh119_16_32 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_16_33 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_16_16 :  std_logic_vector(2 downto 0);
signal heap_bh119_w44_4, heap_bh119_w44_4_d1, heap_bh119_w44_4_d2 :  std_logic;
signal heap_bh119_w45_3, heap_bh119_w45_3_d1, heap_bh119_w45_3_d2 :  std_logic;
signal heap_bh119_w46_3, heap_bh119_w46_3_d1, heap_bh119_w46_3_d2 :  std_logic;
signal CompressorIn_bh119_17_34 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_17_35 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_17_17 :  std_logic_vector(2 downto 0);
signal heap_bh119_w46_4, heap_bh119_w46_4_d1, heap_bh119_w46_4_d2 :  std_logic;
signal heap_bh119_w47_3, heap_bh119_w47_3_d1, heap_bh119_w47_3_d2 :  std_logic;
signal heap_bh119_w48_3, heap_bh119_w48_3_d1, heap_bh119_w48_3_d2 :  std_logic;
signal CompressorIn_bh119_18_36 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_18_37 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_18_18 :  std_logic_vector(2 downto 0);
signal heap_bh119_w48_4, heap_bh119_w48_4_d1, heap_bh119_w48_4_d2 :  std_logic;
signal heap_bh119_w49_3, heap_bh119_w49_3_d1, heap_bh119_w49_3_d2 :  std_logic;
signal heap_bh119_w50_3, heap_bh119_w50_3_d1, heap_bh119_w50_3_d2 :  std_logic;
signal CompressorIn_bh119_19_38 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_19_39 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_19_19 :  std_logic_vector(2 downto 0);
signal heap_bh119_w50_4, heap_bh119_w50_4_d1, heap_bh119_w50_4_d2 :  std_logic;
signal heap_bh119_w51_3, heap_bh119_w51_3_d1, heap_bh119_w51_3_d2 :  std_logic;
signal heap_bh119_w52_3, heap_bh119_w52_3_d1, heap_bh119_w52_3_d2 :  std_logic;
signal CompressorIn_bh119_20_40 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_20_41 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_20_20 :  std_logic_vector(2 downto 0);
signal heap_bh119_w52_4, heap_bh119_w52_4_d1, heap_bh119_w52_4_d2 :  std_logic;
signal heap_bh119_w53_3, heap_bh119_w53_3_d1, heap_bh119_w53_3_d2 :  std_logic;
signal heap_bh119_w54_3, heap_bh119_w54_3_d1, heap_bh119_w54_3_d2 :  std_logic;
signal CompressorIn_bh119_21_42 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_21_43 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_21_21 :  std_logic_vector(2 downto 0);
signal heap_bh119_w54_4, heap_bh119_w54_4_d1, heap_bh119_w54_4_d2 :  std_logic;
signal heap_bh119_w55_3, heap_bh119_w55_3_d1, heap_bh119_w55_3_d2 :  std_logic;
signal heap_bh119_w56_2 :  std_logic;
signal CompressorIn_bh119_22_44 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_22_45 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_22_22 :  std_logic_vector(2 downto 0);
signal heap_bh119_w56_3, heap_bh119_w56_3_d1, heap_bh119_w56_3_d2 :  std_logic;
signal heap_bh119_w57_2, heap_bh119_w57_2_d1, heap_bh119_w57_2_d2 :  std_logic;
signal heap_bh119_w58_2, heap_bh119_w58_2_d1 :  std_logic;
signal CompressorIn_bh119_23_46 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_23_47 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_23_23 :  std_logic_vector(2 downto 0);
signal heap_bh119_w58_3, heap_bh119_w58_3_d1 :  std_logic;
signal heap_bh119_w59_2, heap_bh119_w59_2_d1 :  std_logic;
signal heap_bh119_w60_2 :  std_logic;
signal CompressorIn_bh119_24_48 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh119_24_49 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh119_24_24 :  std_logic_vector(2 downto 0);
signal heap_bh119_w60_3, heap_bh119_w60_3_d1 :  std_logic;
signal heap_bh119_w61_2, heap_bh119_w61_2_d1 :  std_logic;
signal heap_bh119_w62_1, heap_bh119_w62_1_d1 :  std_logic;
signal finalAdderIn0_bh119 :  std_logic_vector(60 downto 0);
signal finalAdderIn1_bh119 :  std_logic_vector(60 downto 0);
signal finalAdderCin_bh119 :  std_logic;
signal finalAdderOut_bh119 :  std_logic_vector(60 downto 0);
signal CompressionResult119 :  std_logic_vector(66 downto 0);
signal OutRes :  std_logic_vector(65 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of KCMTable_4_780414346020670_unsigned_F400_uid112: component is "yes";
attribute rom_extract of KCMTable_6_780414346020670_unsigned_F400_uid110: component is "yes";
attribute rom_style of KCMTable_4_780414346020670_unsigned_F400_uid112: component is "distributed";
attribute rom_style of KCMTable_6_780414346020670_unsigned_F400_uid110: component is "distributed";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            heap_bh119_w6_0_d1 <=  heap_bh119_w6_0;
            heap_bh119_w6_0_d2 <=  heap_bh119_w6_0_d1;
            heap_bh119_w7_0_d1 <=  heap_bh119_w7_0;
            heap_bh119_w7_0_d2 <=  heap_bh119_w7_0_d1;
            heap_bh119_w8_0_d1 <=  heap_bh119_w8_0;
            heap_bh119_w8_0_d2 <=  heap_bh119_w8_0_d1;
            heap_bh119_w9_0_d1 <=  heap_bh119_w9_0;
            heap_bh119_w9_0_d2 <=  heap_bh119_w9_0_d1;
            heap_bh119_w10_0_d1 <=  heap_bh119_w10_0;
            heap_bh119_w10_0_d2 <=  heap_bh119_w10_0_d1;
            heap_bh119_w11_0_d1 <=  heap_bh119_w11_0;
            heap_bh119_w11_0_d2 <=  heap_bh119_w11_0_d1;
            heap_bh119_w13_0_d1 <=  heap_bh119_w13_0;
            heap_bh119_w13_0_d2 <=  heap_bh119_w13_0_d1;
            heap_bh119_w15_0_d1 <=  heap_bh119_w15_0;
            heap_bh119_w15_0_d2 <=  heap_bh119_w15_0_d1;
            heap_bh119_w17_0_d1 <=  heap_bh119_w17_0;
            heap_bh119_w17_0_d2 <=  heap_bh119_w17_0_d1;
            heap_bh119_w19_0_d1 <=  heap_bh119_w19_0;
            heap_bh119_w19_0_d2 <=  heap_bh119_w19_0_d1;
            heap_bh119_w21_0_d1 <=  heap_bh119_w21_0;
            heap_bh119_w21_0_d2 <=  heap_bh119_w21_0_d1;
            heap_bh119_w23_0_d1 <=  heap_bh119_w23_0;
            heap_bh119_w23_0_d2 <=  heap_bh119_w23_0_d1;
            heap_bh119_w25_0_d1 <=  heap_bh119_w25_0;
            heap_bh119_w25_0_d2 <=  heap_bh119_w25_0_d1;
            heap_bh119_w27_0_d1 <=  heap_bh119_w27_0;
            heap_bh119_w27_0_d2 <=  heap_bh119_w27_0_d1;
            heap_bh119_w29_0_d1 <=  heap_bh119_w29_0;
            heap_bh119_w29_0_d2 <=  heap_bh119_w29_0_d1;
            heap_bh119_w31_0_d1 <=  heap_bh119_w31_0;
            heap_bh119_w31_0_d2 <=  heap_bh119_w31_0_d1;
            heap_bh119_w33_0_d1 <=  heap_bh119_w33_0;
            heap_bh119_w33_0_d2 <=  heap_bh119_w33_0_d1;
            heap_bh119_w35_0_d1 <=  heap_bh119_w35_0;
            heap_bh119_w35_0_d2 <=  heap_bh119_w35_0_d1;
            heap_bh119_w37_0_d1 <=  heap_bh119_w37_0;
            heap_bh119_w37_0_d2 <=  heap_bh119_w37_0_d1;
            heap_bh119_w39_0_d1 <=  heap_bh119_w39_0;
            heap_bh119_w39_0_d2 <=  heap_bh119_w39_0_d1;
            heap_bh119_w41_0_d1 <=  heap_bh119_w41_0;
            heap_bh119_w41_0_d2 <=  heap_bh119_w41_0_d1;
            heap_bh119_w43_0_d1 <=  heap_bh119_w43_0;
            heap_bh119_w43_0_d2 <=  heap_bh119_w43_0_d1;
            heap_bh119_w45_0_d1 <=  heap_bh119_w45_0;
            heap_bh119_w45_0_d2 <=  heap_bh119_w45_0_d1;
            heap_bh119_w47_0_d1 <=  heap_bh119_w47_0;
            heap_bh119_w47_0_d2 <=  heap_bh119_w47_0_d1;
            heap_bh119_w49_0_d1 <=  heap_bh119_w49_0;
            heap_bh119_w49_0_d2 <=  heap_bh119_w49_0_d1;
            heap_bh119_w51_0_d1 <=  heap_bh119_w51_0;
            heap_bh119_w51_0_d2 <=  heap_bh119_w51_0_d1;
            heap_bh119_w53_0_d1 <=  heap_bh119_w53_0;
            heap_bh119_w53_0_d2 <=  heap_bh119_w53_0_d1;
            heap_bh119_w55_0_d1 <=  heap_bh119_w55_0;
            heap_bh119_w55_0_d2 <=  heap_bh119_w55_0_d1;
            heap_bh119_w6_1_d1 <=  heap_bh119_w6_1;
            heap_bh119_w6_1_d2 <=  heap_bh119_w6_1_d1;
            heap_bh119_w7_1_d1 <=  heap_bh119_w7_1;
            heap_bh119_w7_1_d2 <=  heap_bh119_w7_1_d1;
            heap_bh119_w8_1_d1 <=  heap_bh119_w8_1;
            heap_bh119_w8_1_d2 <=  heap_bh119_w8_1_d1;
            heap_bh119_w9_1_d1 <=  heap_bh119_w9_1;
            heap_bh119_w9_1_d2 <=  heap_bh119_w9_1_d1;
            heap_bh119_w10_1_d1 <=  heap_bh119_w10_1;
            heap_bh119_w10_1_d2 <=  heap_bh119_w10_1_d1;
            heap_bh119_w11_1_d1 <=  heap_bh119_w11_1;
            heap_bh119_w11_1_d2 <=  heap_bh119_w11_1_d1;
            heap_bh119_w58_0_d1 <=  heap_bh119_w58_0;
            heap_bh119_w59_0_d1 <=  heap_bh119_w59_0;
            heap_bh119_w60_0_d1 <=  heap_bh119_w60_0;
            heap_bh119_w61_0_d1 <=  heap_bh119_w61_0;
            heap_bh119_w58_1_d1 <=  heap_bh119_w58_1;
            heap_bh119_w59_1_d1 <=  heap_bh119_w59_1;
            heap_bh119_w60_1_d1 <=  heap_bh119_w60_1;
            heap_bh119_w61_1_d1 <=  heap_bh119_w61_1;
            heap_bh119_w62_0_d1 <=  heap_bh119_w62_0;
            heap_bh119_w62_0_d2 <=  heap_bh119_w62_0_d1;
            heap_bh119_w63_0_d1 <=  heap_bh119_w63_0;
            heap_bh119_w63_0_d2 <=  heap_bh119_w63_0_d1;
            heap_bh119_w64_0_d1 <=  heap_bh119_w64_0;
            heap_bh119_w64_0_d2 <=  heap_bh119_w64_0_d1;
            heap_bh119_w65_0_d1 <=  heap_bh119_w65_0;
            heap_bh119_w65_0_d2 <=  heap_bh119_w65_0_d1;
            tempR_bh119_0_d1 <=  tempR_bh119_0;
            tempR_bh119_0_d2 <=  tempR_bh119_0_d1;
            tempR_bh119_0_d3 <=  tempR_bh119_0_d2;
            heap_bh119_w12_3_d1 <=  heap_bh119_w12_3;
            heap_bh119_w12_3_d2 <=  heap_bh119_w12_3_d1;
            heap_bh119_w13_3_d1 <=  heap_bh119_w13_3;
            heap_bh119_w13_3_d2 <=  heap_bh119_w13_3_d1;
            heap_bh119_w14_3_d1 <=  heap_bh119_w14_3;
            heap_bh119_w14_3_d2 <=  heap_bh119_w14_3_d1;
            heap_bh119_w14_4_d1 <=  heap_bh119_w14_4;
            heap_bh119_w14_4_d2 <=  heap_bh119_w14_4_d1;
            heap_bh119_w15_3_d1 <=  heap_bh119_w15_3;
            heap_bh119_w15_3_d2 <=  heap_bh119_w15_3_d1;
            heap_bh119_w16_3_d1 <=  heap_bh119_w16_3;
            heap_bh119_w16_3_d2 <=  heap_bh119_w16_3_d1;
            heap_bh119_w16_4_d1 <=  heap_bh119_w16_4;
            heap_bh119_w16_4_d2 <=  heap_bh119_w16_4_d1;
            heap_bh119_w17_3_d1 <=  heap_bh119_w17_3;
            heap_bh119_w17_3_d2 <=  heap_bh119_w17_3_d1;
            heap_bh119_w18_3_d1 <=  heap_bh119_w18_3;
            heap_bh119_w18_3_d2 <=  heap_bh119_w18_3_d1;
            heap_bh119_w18_4_d1 <=  heap_bh119_w18_4;
            heap_bh119_w18_4_d2 <=  heap_bh119_w18_4_d1;
            heap_bh119_w19_3_d1 <=  heap_bh119_w19_3;
            heap_bh119_w19_3_d2 <=  heap_bh119_w19_3_d1;
            heap_bh119_w20_3_d1 <=  heap_bh119_w20_3;
            heap_bh119_w20_3_d2 <=  heap_bh119_w20_3_d1;
            heap_bh119_w20_4_d1 <=  heap_bh119_w20_4;
            heap_bh119_w20_4_d2 <=  heap_bh119_w20_4_d1;
            heap_bh119_w21_3_d1 <=  heap_bh119_w21_3;
            heap_bh119_w21_3_d2 <=  heap_bh119_w21_3_d1;
            heap_bh119_w22_3_d1 <=  heap_bh119_w22_3;
            heap_bh119_w22_3_d2 <=  heap_bh119_w22_3_d1;
            heap_bh119_w22_4_d1 <=  heap_bh119_w22_4;
            heap_bh119_w22_4_d2 <=  heap_bh119_w22_4_d1;
            heap_bh119_w23_3_d1 <=  heap_bh119_w23_3;
            heap_bh119_w23_3_d2 <=  heap_bh119_w23_3_d1;
            heap_bh119_w24_3_d1 <=  heap_bh119_w24_3;
            heap_bh119_w24_3_d2 <=  heap_bh119_w24_3_d1;
            heap_bh119_w24_4_d1 <=  heap_bh119_w24_4;
            heap_bh119_w24_4_d2 <=  heap_bh119_w24_4_d1;
            heap_bh119_w25_3_d1 <=  heap_bh119_w25_3;
            heap_bh119_w25_3_d2 <=  heap_bh119_w25_3_d1;
            heap_bh119_w26_3_d1 <=  heap_bh119_w26_3;
            heap_bh119_w26_3_d2 <=  heap_bh119_w26_3_d1;
            heap_bh119_w26_4_d1 <=  heap_bh119_w26_4;
            heap_bh119_w26_4_d2 <=  heap_bh119_w26_4_d1;
            heap_bh119_w27_3_d1 <=  heap_bh119_w27_3;
            heap_bh119_w27_3_d2 <=  heap_bh119_w27_3_d1;
            heap_bh119_w28_3_d1 <=  heap_bh119_w28_3;
            heap_bh119_w28_3_d2 <=  heap_bh119_w28_3_d1;
            heap_bh119_w28_4_d1 <=  heap_bh119_w28_4;
            heap_bh119_w28_4_d2 <=  heap_bh119_w28_4_d1;
            heap_bh119_w29_3_d1 <=  heap_bh119_w29_3;
            heap_bh119_w29_3_d2 <=  heap_bh119_w29_3_d1;
            heap_bh119_w30_3_d1 <=  heap_bh119_w30_3;
            heap_bh119_w30_3_d2 <=  heap_bh119_w30_3_d1;
            heap_bh119_w30_4_d1 <=  heap_bh119_w30_4;
            heap_bh119_w30_4_d2 <=  heap_bh119_w30_4_d1;
            heap_bh119_w31_3_d1 <=  heap_bh119_w31_3;
            heap_bh119_w31_3_d2 <=  heap_bh119_w31_3_d1;
            heap_bh119_w32_3_d1 <=  heap_bh119_w32_3;
            heap_bh119_w32_3_d2 <=  heap_bh119_w32_3_d1;
            heap_bh119_w32_4_d1 <=  heap_bh119_w32_4;
            heap_bh119_w32_4_d2 <=  heap_bh119_w32_4_d1;
            heap_bh119_w33_3_d1 <=  heap_bh119_w33_3;
            heap_bh119_w33_3_d2 <=  heap_bh119_w33_3_d1;
            heap_bh119_w34_3_d1 <=  heap_bh119_w34_3;
            heap_bh119_w34_3_d2 <=  heap_bh119_w34_3_d1;
            heap_bh119_w34_4_d1 <=  heap_bh119_w34_4;
            heap_bh119_w34_4_d2 <=  heap_bh119_w34_4_d1;
            heap_bh119_w35_3_d1 <=  heap_bh119_w35_3;
            heap_bh119_w35_3_d2 <=  heap_bh119_w35_3_d1;
            heap_bh119_w36_3_d1 <=  heap_bh119_w36_3;
            heap_bh119_w36_3_d2 <=  heap_bh119_w36_3_d1;
            heap_bh119_w36_4_d1 <=  heap_bh119_w36_4;
            heap_bh119_w36_4_d2 <=  heap_bh119_w36_4_d1;
            heap_bh119_w37_3_d1 <=  heap_bh119_w37_3;
            heap_bh119_w37_3_d2 <=  heap_bh119_w37_3_d1;
            heap_bh119_w38_3_d1 <=  heap_bh119_w38_3;
            heap_bh119_w38_3_d2 <=  heap_bh119_w38_3_d1;
            heap_bh119_w38_4_d1 <=  heap_bh119_w38_4;
            heap_bh119_w38_4_d2 <=  heap_bh119_w38_4_d1;
            heap_bh119_w39_3_d1 <=  heap_bh119_w39_3;
            heap_bh119_w39_3_d2 <=  heap_bh119_w39_3_d1;
            heap_bh119_w40_3_d1 <=  heap_bh119_w40_3;
            heap_bh119_w40_3_d2 <=  heap_bh119_w40_3_d1;
            heap_bh119_w40_4_d1 <=  heap_bh119_w40_4;
            heap_bh119_w40_4_d2 <=  heap_bh119_w40_4_d1;
            heap_bh119_w41_3_d1 <=  heap_bh119_w41_3;
            heap_bh119_w41_3_d2 <=  heap_bh119_w41_3_d1;
            heap_bh119_w42_3_d1 <=  heap_bh119_w42_3;
            heap_bh119_w42_3_d2 <=  heap_bh119_w42_3_d1;
            heap_bh119_w42_4_d1 <=  heap_bh119_w42_4;
            heap_bh119_w42_4_d2 <=  heap_bh119_w42_4_d1;
            heap_bh119_w43_3_d1 <=  heap_bh119_w43_3;
            heap_bh119_w43_3_d2 <=  heap_bh119_w43_3_d1;
            heap_bh119_w44_3_d1 <=  heap_bh119_w44_3;
            heap_bh119_w44_3_d2 <=  heap_bh119_w44_3_d1;
            heap_bh119_w44_4_d1 <=  heap_bh119_w44_4;
            heap_bh119_w44_4_d2 <=  heap_bh119_w44_4_d1;
            heap_bh119_w45_3_d1 <=  heap_bh119_w45_3;
            heap_bh119_w45_3_d2 <=  heap_bh119_w45_3_d1;
            heap_bh119_w46_3_d1 <=  heap_bh119_w46_3;
            heap_bh119_w46_3_d2 <=  heap_bh119_w46_3_d1;
            heap_bh119_w46_4_d1 <=  heap_bh119_w46_4;
            heap_bh119_w46_4_d2 <=  heap_bh119_w46_4_d1;
            heap_bh119_w47_3_d1 <=  heap_bh119_w47_3;
            heap_bh119_w47_3_d2 <=  heap_bh119_w47_3_d1;
            heap_bh119_w48_3_d1 <=  heap_bh119_w48_3;
            heap_bh119_w48_3_d2 <=  heap_bh119_w48_3_d1;
            heap_bh119_w48_4_d1 <=  heap_bh119_w48_4;
            heap_bh119_w48_4_d2 <=  heap_bh119_w48_4_d1;
            heap_bh119_w49_3_d1 <=  heap_bh119_w49_3;
            heap_bh119_w49_3_d2 <=  heap_bh119_w49_3_d1;
            heap_bh119_w50_3_d1 <=  heap_bh119_w50_3;
            heap_bh119_w50_3_d2 <=  heap_bh119_w50_3_d1;
            heap_bh119_w50_4_d1 <=  heap_bh119_w50_4;
            heap_bh119_w50_4_d2 <=  heap_bh119_w50_4_d1;
            heap_bh119_w51_3_d1 <=  heap_bh119_w51_3;
            heap_bh119_w51_3_d2 <=  heap_bh119_w51_3_d1;
            heap_bh119_w52_3_d1 <=  heap_bh119_w52_3;
            heap_bh119_w52_3_d2 <=  heap_bh119_w52_3_d1;
            heap_bh119_w52_4_d1 <=  heap_bh119_w52_4;
            heap_bh119_w52_4_d2 <=  heap_bh119_w52_4_d1;
            heap_bh119_w53_3_d1 <=  heap_bh119_w53_3;
            heap_bh119_w53_3_d2 <=  heap_bh119_w53_3_d1;
            heap_bh119_w54_3_d1 <=  heap_bh119_w54_3;
            heap_bh119_w54_3_d2 <=  heap_bh119_w54_3_d1;
            heap_bh119_w54_4_d1 <=  heap_bh119_w54_4;
            heap_bh119_w54_4_d2 <=  heap_bh119_w54_4_d1;
            heap_bh119_w55_3_d1 <=  heap_bh119_w55_3;
            heap_bh119_w55_3_d2 <=  heap_bh119_w55_3_d1;
            heap_bh119_w56_3_d1 <=  heap_bh119_w56_3;
            heap_bh119_w56_3_d2 <=  heap_bh119_w56_3_d1;
            heap_bh119_w57_2_d1 <=  heap_bh119_w57_2;
            heap_bh119_w57_2_d2 <=  heap_bh119_w57_2_d1;
            heap_bh119_w58_2_d1 <=  heap_bh119_w58_2;
            heap_bh119_w58_3_d1 <=  heap_bh119_w58_3;
            heap_bh119_w59_2_d1 <=  heap_bh119_w59_2;
            heap_bh119_w60_3_d1 <=  heap_bh119_w60_3;
            heap_bh119_w61_2_d1 <=  heap_bh119_w61_2;
            heap_bh119_w62_1_d1 <=  heap_bh119_w62_1;
         end if;
      end process;
   d0 <= X(5 downto 0);
   KCMTable_0: KCMTable_6_780414346020670_unsigned_F400_uid110  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => d0,
                 Y => pp0);
   d1 <= X(11 downto 6);
   KCMTable_1: KCMTable_6_780414346020670_unsigned_F400_uid110  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => d1,
                 Y => pp1);
   d2 <= X(15 downto 12);
   KCMTable_2: KCMTable_4_780414346020670_unsigned_F400_uid112  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => d2,
                 Y => pp2);
   heap_bh119_w0_0 <= pp0(0); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w1_0 <= pp0(1); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w2_0 <= pp0(2); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w3_0 <= pp0(3); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w4_0 <= pp0(4); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w5_0 <= pp0(5); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w6_0 <= pp0(6); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w7_0 <= pp0(7); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w8_0 <= pp0(8); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w9_0 <= pp0(9); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w10_0 <= pp0(10); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w11_0 <= pp0(11); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w12_0 <= pp0(12); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w13_0 <= pp0(13); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w14_0 <= pp0(14); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w15_0 <= pp0(15); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w16_0 <= pp0(16); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w17_0 <= pp0(17); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w18_0 <= pp0(18); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w19_0 <= pp0(19); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w20_0 <= pp0(20); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w21_0 <= pp0(21); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w22_0 <= pp0(22); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w23_0 <= pp0(23); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w24_0 <= pp0(24); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w25_0 <= pp0(25); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w26_0 <= pp0(26); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w27_0 <= pp0(27); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w28_0 <= pp0(28); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w29_0 <= pp0(29); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w30_0 <= pp0(30); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w31_0 <= pp0(31); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w32_0 <= pp0(32); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w33_0 <= pp0(33); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w34_0 <= pp0(34); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w35_0 <= pp0(35); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w36_0 <= pp0(36); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w37_0 <= pp0(37); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w38_0 <= pp0(38); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w39_0 <= pp0(39); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w40_0 <= pp0(40); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w41_0 <= pp0(41); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w42_0 <= pp0(42); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w43_0 <= pp0(43); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w44_0 <= pp0(44); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w45_0 <= pp0(45); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w46_0 <= pp0(46); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w47_0 <= pp0(47); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w48_0 <= pp0(48); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w49_0 <= pp0(49); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w50_0 <= pp0(50); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w51_0 <= pp0(51); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w52_0 <= pp0(52); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w53_0 <= pp0(53); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w54_0 <= pp0(54); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w55_0 <= pp0(55); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w6_1 <= pp1(0); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w7_1 <= pp1(1); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w8_1 <= pp1(2); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w9_1 <= pp1(3); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w10_1 <= pp1(4); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w11_1 <= pp1(5); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w12_1 <= pp1(6); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w13_1 <= pp1(7); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w14_1 <= pp1(8); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w15_1 <= pp1(9); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w16_1 <= pp1(10); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w17_1 <= pp1(11); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w18_1 <= pp1(12); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w19_1 <= pp1(13); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w20_1 <= pp1(14); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w21_1 <= pp1(15); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w22_1 <= pp1(16); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w23_1 <= pp1(17); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w24_1 <= pp1(18); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w25_1 <= pp1(19); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w26_1 <= pp1(20); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w27_1 <= pp1(21); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w28_1 <= pp1(22); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w29_1 <= pp1(23); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w30_1 <= pp1(24); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w31_1 <= pp1(25); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w32_1 <= pp1(26); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w33_1 <= pp1(27); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w34_1 <= pp1(28); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w35_1 <= pp1(29); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w36_1 <= pp1(30); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w37_1 <= pp1(31); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w38_1 <= pp1(32); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w39_1 <= pp1(33); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w40_1 <= pp1(34); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w41_1 <= pp1(35); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w42_1 <= pp1(36); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w43_1 <= pp1(37); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w44_1 <= pp1(38); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w45_1 <= pp1(39); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w46_1 <= pp1(40); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w47_1 <= pp1(41); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w48_1 <= pp1(42); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w49_1 <= pp1(43); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w50_1 <= pp1(44); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w51_1 <= pp1(45); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w52_1 <= pp1(46); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w53_1 <= pp1(47); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w54_1 <= pp1(48); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w55_1 <= pp1(49); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w56_0 <= pp1(50); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w57_0 <= pp1(51); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w58_0 <= pp1(52); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w59_0 <= pp1(53); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w60_0 <= pp1(54); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w61_0 <= pp1(55); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w12_2 <= pp2(0); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w13_2 <= pp2(1); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w14_2 <= pp2(2); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w15_2 <= pp2(3); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w16_2 <= pp2(4); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w17_2 <= pp2(5); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w18_2 <= pp2(6); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w19_2 <= pp2(7); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w20_2 <= pp2(8); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w21_2 <= pp2(9); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w22_2 <= pp2(10); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w23_2 <= pp2(11); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w24_2 <= pp2(12); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w25_2 <= pp2(13); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w26_2 <= pp2(14); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w27_2 <= pp2(15); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w28_2 <= pp2(16); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w29_2 <= pp2(17); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w30_2 <= pp2(18); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w31_2 <= pp2(19); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w32_2 <= pp2(20); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w33_2 <= pp2(21); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w34_2 <= pp2(22); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w35_2 <= pp2(23); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w36_2 <= pp2(24); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w37_2 <= pp2(25); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w38_2 <= pp2(26); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w39_2 <= pp2(27); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w40_2 <= pp2(28); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w41_2 <= pp2(29); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w42_2 <= pp2(30); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w43_2 <= pp2(31); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w44_2 <= pp2(32); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w45_2 <= pp2(33); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w46_2 <= pp2(34); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w47_2 <= pp2(35); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w48_2 <= pp2(36); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w49_2 <= pp2(37); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w50_2 <= pp2(38); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w51_2 <= pp2(39); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w52_2 <= pp2(40); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w53_2 <= pp2(41); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w54_2 <= pp2(42); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w55_2 <= pp2(43); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w56_1 <= pp2(44); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w57_1 <= pp2(45); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w58_1 <= pp2(46); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w59_1 <= pp2(47); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w60_1 <= pp2(48); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w61_1 <= pp2(49); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w62_0 <= pp2(50); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w63_0 <= pp2(51); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w64_0 <= pp2(52); -- cycle= 0 cp= 9.9288e-10
   heap_bh119_w65_0 <= pp2(53); -- cycle= 0 cp= 9.9288e-10
   
   -- Beginning of code generated by BitHeap::generateCompressorVHDL
   -- code generated by BitHeap::generateSupertileVHDL()
   ----------------Synchro barrier, entering cycle 0----------------

   -- Adding the constant bits
      -- All the constant bits are zero, nothing to add

   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 0----------------
   tempR_bh119_0 <= heap_bh119_w5_0 & heap_bh119_w4_0 & heap_bh119_w3_0 & heap_bh119_w2_0 & heap_bh119_w1_0 & heap_bh119_w0_0; -- already compressed

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_0_0 <= heap_bh119_w12_2 & heap_bh119_w12_1 & heap_bh119_w12_0;
   CompressorIn_bh119_0_1 <= heap_bh119_w13_2 & heap_bh119_w13_1;
   Compressor_bh119_0: Compressor_23_3
      port map ( R => CompressorOut_bh119_0_0   ,
                 X0 => CompressorIn_bh119_0_0,
                 X1 => CompressorIn_bh119_0_1);
   heap_bh119_w12_3 <= CompressorOut_bh119_0_0(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w13_3 <= CompressorOut_bh119_0_0(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w14_3 <= CompressorOut_bh119_0_0(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_1_2 <= heap_bh119_w14_2 & heap_bh119_w14_1 & heap_bh119_w14_0;
   CompressorIn_bh119_1_3 <= heap_bh119_w15_2 & heap_bh119_w15_1;
   Compressor_bh119_1: Compressor_23_3
      port map ( R => CompressorOut_bh119_1_1   ,
                 X0 => CompressorIn_bh119_1_2,
                 X1 => CompressorIn_bh119_1_3);
   heap_bh119_w14_4 <= CompressorOut_bh119_1_1(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w15_3 <= CompressorOut_bh119_1_1(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w16_3 <= CompressorOut_bh119_1_1(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_2_4 <= heap_bh119_w16_2 & heap_bh119_w16_1 & heap_bh119_w16_0;
   CompressorIn_bh119_2_5 <= heap_bh119_w17_2 & heap_bh119_w17_1;
   Compressor_bh119_2: Compressor_23_3
      port map ( R => CompressorOut_bh119_2_2   ,
                 X0 => CompressorIn_bh119_2_4,
                 X1 => CompressorIn_bh119_2_5);
   heap_bh119_w16_4 <= CompressorOut_bh119_2_2(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w17_3 <= CompressorOut_bh119_2_2(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w18_3 <= CompressorOut_bh119_2_2(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_3_6 <= heap_bh119_w18_2 & heap_bh119_w18_1 & heap_bh119_w18_0;
   CompressorIn_bh119_3_7 <= heap_bh119_w19_2 & heap_bh119_w19_1;
   Compressor_bh119_3: Compressor_23_3
      port map ( R => CompressorOut_bh119_3_3   ,
                 X0 => CompressorIn_bh119_3_6,
                 X1 => CompressorIn_bh119_3_7);
   heap_bh119_w18_4 <= CompressorOut_bh119_3_3(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w19_3 <= CompressorOut_bh119_3_3(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w20_3 <= CompressorOut_bh119_3_3(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_4_8 <= heap_bh119_w20_2 & heap_bh119_w20_1 & heap_bh119_w20_0;
   CompressorIn_bh119_4_9 <= heap_bh119_w21_2 & heap_bh119_w21_1;
   Compressor_bh119_4: Compressor_23_3
      port map ( R => CompressorOut_bh119_4_4   ,
                 X0 => CompressorIn_bh119_4_8,
                 X1 => CompressorIn_bh119_4_9);
   heap_bh119_w20_4 <= CompressorOut_bh119_4_4(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w21_3 <= CompressorOut_bh119_4_4(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w22_3 <= CompressorOut_bh119_4_4(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_5_10 <= heap_bh119_w22_2 & heap_bh119_w22_1 & heap_bh119_w22_0;
   CompressorIn_bh119_5_11 <= heap_bh119_w23_2 & heap_bh119_w23_1;
   Compressor_bh119_5: Compressor_23_3
      port map ( R => CompressorOut_bh119_5_5   ,
                 X0 => CompressorIn_bh119_5_10,
                 X1 => CompressorIn_bh119_5_11);
   heap_bh119_w22_4 <= CompressorOut_bh119_5_5(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w23_3 <= CompressorOut_bh119_5_5(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w24_3 <= CompressorOut_bh119_5_5(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_6_12 <= heap_bh119_w24_2 & heap_bh119_w24_1 & heap_bh119_w24_0;
   CompressorIn_bh119_6_13 <= heap_bh119_w25_2 & heap_bh119_w25_1;
   Compressor_bh119_6: Compressor_23_3
      port map ( R => CompressorOut_bh119_6_6   ,
                 X0 => CompressorIn_bh119_6_12,
                 X1 => CompressorIn_bh119_6_13);
   heap_bh119_w24_4 <= CompressorOut_bh119_6_6(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w25_3 <= CompressorOut_bh119_6_6(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w26_3 <= CompressorOut_bh119_6_6(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_7_14 <= heap_bh119_w26_2 & heap_bh119_w26_1 & heap_bh119_w26_0;
   CompressorIn_bh119_7_15 <= heap_bh119_w27_2 & heap_bh119_w27_1;
   Compressor_bh119_7: Compressor_23_3
      port map ( R => CompressorOut_bh119_7_7   ,
                 X0 => CompressorIn_bh119_7_14,
                 X1 => CompressorIn_bh119_7_15);
   heap_bh119_w26_4 <= CompressorOut_bh119_7_7(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w27_3 <= CompressorOut_bh119_7_7(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w28_3 <= CompressorOut_bh119_7_7(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_8_16 <= heap_bh119_w28_2 & heap_bh119_w28_1 & heap_bh119_w28_0;
   CompressorIn_bh119_8_17 <= heap_bh119_w29_2 & heap_bh119_w29_1;
   Compressor_bh119_8: Compressor_23_3
      port map ( R => CompressorOut_bh119_8_8   ,
                 X0 => CompressorIn_bh119_8_16,
                 X1 => CompressorIn_bh119_8_17);
   heap_bh119_w28_4 <= CompressorOut_bh119_8_8(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w29_3 <= CompressorOut_bh119_8_8(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w30_3 <= CompressorOut_bh119_8_8(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_9_18 <= heap_bh119_w30_2 & heap_bh119_w30_1 & heap_bh119_w30_0;
   CompressorIn_bh119_9_19 <= heap_bh119_w31_2 & heap_bh119_w31_1;
   Compressor_bh119_9: Compressor_23_3
      port map ( R => CompressorOut_bh119_9_9   ,
                 X0 => CompressorIn_bh119_9_18,
                 X1 => CompressorIn_bh119_9_19);
   heap_bh119_w30_4 <= CompressorOut_bh119_9_9(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w31_3 <= CompressorOut_bh119_9_9(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w32_3 <= CompressorOut_bh119_9_9(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_10_20 <= heap_bh119_w32_2 & heap_bh119_w32_1 & heap_bh119_w32_0;
   CompressorIn_bh119_10_21 <= heap_bh119_w33_2 & heap_bh119_w33_1;
   Compressor_bh119_10: Compressor_23_3
      port map ( R => CompressorOut_bh119_10_10   ,
                 X0 => CompressorIn_bh119_10_20,
                 X1 => CompressorIn_bh119_10_21);
   heap_bh119_w32_4 <= CompressorOut_bh119_10_10(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w33_3 <= CompressorOut_bh119_10_10(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w34_3 <= CompressorOut_bh119_10_10(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_11_22 <= heap_bh119_w34_2 & heap_bh119_w34_1 & heap_bh119_w34_0;
   CompressorIn_bh119_11_23 <= heap_bh119_w35_2 & heap_bh119_w35_1;
   Compressor_bh119_11: Compressor_23_3
      port map ( R => CompressorOut_bh119_11_11   ,
                 X0 => CompressorIn_bh119_11_22,
                 X1 => CompressorIn_bh119_11_23);
   heap_bh119_w34_4 <= CompressorOut_bh119_11_11(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w35_3 <= CompressorOut_bh119_11_11(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w36_3 <= CompressorOut_bh119_11_11(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_12_24 <= heap_bh119_w36_2 & heap_bh119_w36_1 & heap_bh119_w36_0;
   CompressorIn_bh119_12_25 <= heap_bh119_w37_2 & heap_bh119_w37_1;
   Compressor_bh119_12: Compressor_23_3
      port map ( R => CompressorOut_bh119_12_12   ,
                 X0 => CompressorIn_bh119_12_24,
                 X1 => CompressorIn_bh119_12_25);
   heap_bh119_w36_4 <= CompressorOut_bh119_12_12(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w37_3 <= CompressorOut_bh119_12_12(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w38_3 <= CompressorOut_bh119_12_12(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_13_26 <= heap_bh119_w38_2 & heap_bh119_w38_1 & heap_bh119_w38_0;
   CompressorIn_bh119_13_27 <= heap_bh119_w39_2 & heap_bh119_w39_1;
   Compressor_bh119_13: Compressor_23_3
      port map ( R => CompressorOut_bh119_13_13   ,
                 X0 => CompressorIn_bh119_13_26,
                 X1 => CompressorIn_bh119_13_27);
   heap_bh119_w38_4 <= CompressorOut_bh119_13_13(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w39_3 <= CompressorOut_bh119_13_13(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w40_3 <= CompressorOut_bh119_13_13(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_14_28 <= heap_bh119_w40_2 & heap_bh119_w40_1 & heap_bh119_w40_0;
   CompressorIn_bh119_14_29 <= heap_bh119_w41_2 & heap_bh119_w41_1;
   Compressor_bh119_14: Compressor_23_3
      port map ( R => CompressorOut_bh119_14_14   ,
                 X0 => CompressorIn_bh119_14_28,
                 X1 => CompressorIn_bh119_14_29);
   heap_bh119_w40_4 <= CompressorOut_bh119_14_14(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w41_3 <= CompressorOut_bh119_14_14(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w42_3 <= CompressorOut_bh119_14_14(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_15_30 <= heap_bh119_w42_2 & heap_bh119_w42_1 & heap_bh119_w42_0;
   CompressorIn_bh119_15_31 <= heap_bh119_w43_2 & heap_bh119_w43_1;
   Compressor_bh119_15: Compressor_23_3
      port map ( R => CompressorOut_bh119_15_15   ,
                 X0 => CompressorIn_bh119_15_30,
                 X1 => CompressorIn_bh119_15_31);
   heap_bh119_w42_4 <= CompressorOut_bh119_15_15(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w43_3 <= CompressorOut_bh119_15_15(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w44_3 <= CompressorOut_bh119_15_15(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_16_32 <= heap_bh119_w44_2 & heap_bh119_w44_1 & heap_bh119_w44_0;
   CompressorIn_bh119_16_33 <= heap_bh119_w45_2 & heap_bh119_w45_1;
   Compressor_bh119_16: Compressor_23_3
      port map ( R => CompressorOut_bh119_16_16   ,
                 X0 => CompressorIn_bh119_16_32,
                 X1 => CompressorIn_bh119_16_33);
   heap_bh119_w44_4 <= CompressorOut_bh119_16_16(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w45_3 <= CompressorOut_bh119_16_16(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w46_3 <= CompressorOut_bh119_16_16(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_17_34 <= heap_bh119_w46_2 & heap_bh119_w46_1 & heap_bh119_w46_0;
   CompressorIn_bh119_17_35 <= heap_bh119_w47_2 & heap_bh119_w47_1;
   Compressor_bh119_17: Compressor_23_3
      port map ( R => CompressorOut_bh119_17_17   ,
                 X0 => CompressorIn_bh119_17_34,
                 X1 => CompressorIn_bh119_17_35);
   heap_bh119_w46_4 <= CompressorOut_bh119_17_17(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w47_3 <= CompressorOut_bh119_17_17(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w48_3 <= CompressorOut_bh119_17_17(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_18_36 <= heap_bh119_w48_2 & heap_bh119_w48_1 & heap_bh119_w48_0;
   CompressorIn_bh119_18_37 <= heap_bh119_w49_2 & heap_bh119_w49_1;
   Compressor_bh119_18: Compressor_23_3
      port map ( R => CompressorOut_bh119_18_18   ,
                 X0 => CompressorIn_bh119_18_36,
                 X1 => CompressorIn_bh119_18_37);
   heap_bh119_w48_4 <= CompressorOut_bh119_18_18(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w49_3 <= CompressorOut_bh119_18_18(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w50_3 <= CompressorOut_bh119_18_18(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_19_38 <= heap_bh119_w50_2 & heap_bh119_w50_1 & heap_bh119_w50_0;
   CompressorIn_bh119_19_39 <= heap_bh119_w51_2 & heap_bh119_w51_1;
   Compressor_bh119_19: Compressor_23_3
      port map ( R => CompressorOut_bh119_19_19   ,
                 X0 => CompressorIn_bh119_19_38,
                 X1 => CompressorIn_bh119_19_39);
   heap_bh119_w50_4 <= CompressorOut_bh119_19_19(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w51_3 <= CompressorOut_bh119_19_19(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w52_3 <= CompressorOut_bh119_19_19(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_20_40 <= heap_bh119_w52_2 & heap_bh119_w52_1 & heap_bh119_w52_0;
   CompressorIn_bh119_20_41 <= heap_bh119_w53_2 & heap_bh119_w53_1;
   Compressor_bh119_20: Compressor_23_3
      port map ( R => CompressorOut_bh119_20_20   ,
                 X0 => CompressorIn_bh119_20_40,
                 X1 => CompressorIn_bh119_20_41);
   heap_bh119_w52_4 <= CompressorOut_bh119_20_20(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w53_3 <= CompressorOut_bh119_20_20(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w54_3 <= CompressorOut_bh119_20_20(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_21_42 <= heap_bh119_w54_2 & heap_bh119_w54_1 & heap_bh119_w54_0;
   CompressorIn_bh119_21_43 <= heap_bh119_w55_2 & heap_bh119_w55_1;
   Compressor_bh119_21: Compressor_23_3
      port map ( R => CompressorOut_bh119_21_21   ,
                 X0 => CompressorIn_bh119_21_42,
                 X1 => CompressorIn_bh119_21_43);
   heap_bh119_w54_4 <= CompressorOut_bh119_21_21(0); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w55_3 <= CompressorOut_bh119_21_21(1); -- cycle= 0 cp= 1.5236e-09
   heap_bh119_w56_2 <= CompressorOut_bh119_21_21(2); -- cycle= 0 cp= 1.5236e-09

   ----------------Synchro barrier, entering cycle 0----------------
   CompressorIn_bh119_22_44 <= heap_bh119_w56_1 & heap_bh119_w56_0 & heap_bh119_w56_2;
   CompressorIn_bh119_22_45 <= heap_bh119_w57_1 & heap_bh119_w57_0;
   Compressor_bh119_22: Compressor_23_3
      port map ( R => CompressorOut_bh119_22_22   ,
                 X0 => CompressorIn_bh119_22_44,
                 X1 => CompressorIn_bh119_22_45);
   heap_bh119_w56_3 <= CompressorOut_bh119_22_22(0); -- cycle= 0 cp= 2.05432e-09
   heap_bh119_w57_2 <= CompressorOut_bh119_22_22(1); -- cycle= 0 cp= 2.05432e-09
   heap_bh119_w58_2 <= CompressorOut_bh119_22_22(2); -- cycle= 0 cp= 2.05432e-09

   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   CompressorIn_bh119_23_46 <= heap_bh119_w58_1_d1 & heap_bh119_w58_0_d1 & heap_bh119_w58_2_d1;
   CompressorIn_bh119_23_47 <= heap_bh119_w59_1_d1 & heap_bh119_w59_0_d1;
   Compressor_bh119_23: Compressor_23_3
      port map ( R => CompressorOut_bh119_23_23   ,
                 X0 => CompressorIn_bh119_23_46,
                 X1 => CompressorIn_bh119_23_47);
   heap_bh119_w58_3 <= CompressorOut_bh119_23_23(0); -- cycle= 1 cp= 0
   heap_bh119_w59_2 <= CompressorOut_bh119_23_23(1); -- cycle= 1 cp= 0
   heap_bh119_w60_2 <= CompressorOut_bh119_23_23(2); -- cycle= 1 cp= 0

   ----------------Synchro barrier, entering cycle 1----------------
   CompressorIn_bh119_24_48 <= heap_bh119_w60_1_d1 & heap_bh119_w60_0_d1 & heap_bh119_w60_2;
   CompressorIn_bh119_24_49 <= heap_bh119_w61_1_d1 & heap_bh119_w61_0_d1;
   Compressor_bh119_24: Compressor_23_3
      port map ( R => CompressorOut_bh119_24_24   ,
                 X0 => CompressorIn_bh119_24_48,
                 X1 => CompressorIn_bh119_24_49);
   heap_bh119_w60_3 <= CompressorOut_bh119_24_24(0); -- cycle= 1 cp= 5.3072e-10
   heap_bh119_w61_2 <= CompressorOut_bh119_24_24(1); -- cycle= 1 cp= 5.3072e-10
   heap_bh119_w62_1 <= CompressorOut_bh119_24_24(2); -- cycle= 1 cp= 5.3072e-10
   ----------------Synchro barrier, entering cycle 1----------------
   ----------------Synchro barrier, entering cycle 2----------------
   finalAdderIn0_bh119 <= "0" & heap_bh119_w65_0_d2 & heap_bh119_w64_0_d2 & heap_bh119_w63_0_d2 & heap_bh119_w62_0_d2 & heap_bh119_w61_2_d1 & heap_bh119_w60_3_d1 & heap_bh119_w59_2_d1 & heap_bh119_w58_3_d1 & heap_bh119_w57_2_d2 & heap_bh119_w56_3_d2 & heap_bh119_w55_0_d2 & heap_bh119_w54_4_d2 & heap_bh119_w53_0_d2 & heap_bh119_w52_4_d2 & heap_bh119_w51_0_d2 & heap_bh119_w50_4_d2 & heap_bh119_w49_0_d2 & heap_bh119_w48_4_d2 & heap_bh119_w47_0_d2 & heap_bh119_w46_4_d2 & heap_bh119_w45_0_d2 & heap_bh119_w44_4_d2 & heap_bh119_w43_0_d2 & heap_bh119_w42_4_d2 & heap_bh119_w41_0_d2 & heap_bh119_w40_4_d2 & heap_bh119_w39_0_d2 & heap_bh119_w38_4_d2 & heap_bh119_w37_0_d2 & heap_bh119_w36_4_d2 & heap_bh119_w35_0_d2 & heap_bh119_w34_4_d2 & heap_bh119_w33_0_d2 & heap_bh119_w32_4_d2 & heap_bh119_w31_0_d2 & heap_bh119_w30_4_d2 & heap_bh119_w29_0_d2 & heap_bh119_w28_4_d2 & heap_bh119_w27_0_d2 & heap_bh119_w26_4_d2 & heap_bh119_w25_0_d2 & heap_bh119_w24_4_d2 & heap_bh119_w23_0_d2 & heap_bh119_w22_4_d2 & heap_bh119_w21_0_d2 & heap_bh119_w20_4_d2 & heap_bh119_w19_0_d2 & heap_bh119_w18_4_d2 & heap_bh119_w17_0_d2 & heap_bh119_w16_4_d2 & heap_bh119_w15_0_d2 & heap_bh119_w14_4_d2 & heap_bh119_w13_0_d2 & heap_bh119_w12_3_d2 & heap_bh119_w11_1_d2 & heap_bh119_w10_1_d2 & heap_bh119_w9_1_d2 & heap_bh119_w8_1_d2 & heap_bh119_w7_1_d2 & heap_bh119_w6_1_d2;
   finalAdderIn1_bh119 <= "0" & '0' & '0' & '0' & heap_bh119_w62_1_d1 & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh119_w55_3_d2 & heap_bh119_w54_3_d2 & heap_bh119_w53_3_d2 & heap_bh119_w52_3_d2 & heap_bh119_w51_3_d2 & heap_bh119_w50_3_d2 & heap_bh119_w49_3_d2 & heap_bh119_w48_3_d2 & heap_bh119_w47_3_d2 & heap_bh119_w46_3_d2 & heap_bh119_w45_3_d2 & heap_bh119_w44_3_d2 & heap_bh119_w43_3_d2 & heap_bh119_w42_3_d2 & heap_bh119_w41_3_d2 & heap_bh119_w40_3_d2 & heap_bh119_w39_3_d2 & heap_bh119_w38_3_d2 & heap_bh119_w37_3_d2 & heap_bh119_w36_3_d2 & heap_bh119_w35_3_d2 & heap_bh119_w34_3_d2 & heap_bh119_w33_3_d2 & heap_bh119_w32_3_d2 & heap_bh119_w31_3_d2 & heap_bh119_w30_3_d2 & heap_bh119_w29_3_d2 & heap_bh119_w28_3_d2 & heap_bh119_w27_3_d2 & heap_bh119_w26_3_d2 & heap_bh119_w25_3_d2 & heap_bh119_w24_3_d2 & heap_bh119_w23_3_d2 & heap_bh119_w22_3_d2 & heap_bh119_w21_3_d2 & heap_bh119_w20_3_d2 & heap_bh119_w19_3_d2 & heap_bh119_w18_3_d2 & heap_bh119_w17_3_d2 & heap_bh119_w16_3_d2 & heap_bh119_w15_3_d2 & heap_bh119_w14_3_d2 & heap_bh119_w13_3_d2 & '0' & heap_bh119_w11_0_d2 & heap_bh119_w10_0_d2 & heap_bh119_w9_0_d2 & heap_bh119_w8_0_d2 & heap_bh119_w7_0_d2 & heap_bh119_w6_0_d2;
   finalAdderCin_bh119 <= '0';
   Adder_final119_0: IntAdder_61_f400_uid178  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => finalAdderCin_bh119,
                 R => finalAdderOut_bh119   ,
                 X => finalAdderIn0_bh119,
                 Y => finalAdderIn1_bh119);
   ----------------Synchro barrier, entering cycle 3----------------
   -- concatenate all the compressed chunks
   CompressionResult119 <= finalAdderOut_bh119 & tempR_bh119_0_d3;
   -- End of code generated by BitHeap::generateCompressorVHDL
OutRes <= CompressionResult119(65 downto 0);
   R <= OutRes;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_90_f400_uid188
--                     (IntAdderClassical_90_F400_uid190)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_90_f400_uid188 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(89 downto 0);
          Y : in  std_logic_vector(89 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(89 downto 0)   );
end entity;

architecture arch of IntAdder_90_f400_uid188 is
signal x0 :  std_logic_vector(13 downto 0);
signal y0 :  std_logic_vector(13 downto 0);
signal x1, x1_d1 :  std_logic_vector(41 downto 0);
signal y1, y1_d1 :  std_logic_vector(41 downto 0);
signal x2, x2_d1, x2_d2 :  std_logic_vector(33 downto 0);
signal y2, y2_d1, y2_d2 :  std_logic_vector(33 downto 0);
signal sum0, sum0_d1, sum0_d2 :  std_logic_vector(14 downto 0);
signal sum1, sum1_d1 :  std_logic_vector(42 downto 0);
signal sum2 :  std_logic_vector(34 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            x1_d1 <=  x1;
            y1_d1 <=  y1;
            x2_d1 <=  x2;
            x2_d2 <=  x2_d1;
            y2_d1 <=  y2;
            y2_d2 <=  y2_d1;
            sum0_d1 <=  sum0;
            sum0_d2 <=  sum0_d1;
            sum1_d1 <=  sum1;
         end if;
      end process;
   --Classical
   x0 <= X(13 downto 0);
   y0 <= Y(13 downto 0);
   x1 <= X(55 downto 14);
   y1 <= Y(55 downto 14);
   x2 <= X(89 downto 56);
   y2 <= Y(89 downto 56);
   sum0 <= ( "0" & x0) + ( "0" & y0)  + Cin;
   ----------------Synchro barrier, entering cycle 1----------------
   sum1 <= ( "0" & x1_d1) + ( "0" & y1_d1)  + sum0_d1(14);
   ----------------Synchro barrier, entering cycle 2----------------
   sum2 <= ( "0" & x2_d2) + ( "0" & y2_d2)  + sum1_d1(42);
   R <= sum2(33 downto 0) & sum1_d1(41 downto 0) & sum0_d2(13 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                LZCShifter_90_to_74_counting_128_F400_uid196
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZCShifter_90_to_74_counting_128_F400_uid196 is
   port ( clk, rst : in std_logic;
          I : in  std_logic_vector(89 downto 0);
          Count : out  std_logic_vector(6 downto 0);
          O : out  std_logic_vector(73 downto 0)   );
end entity;

architecture arch of LZCShifter_90_to_74_counting_128_F400_uid196 is
signal level7, level7_d1 :  std_logic_vector(89 downto 0);
signal count6, count6_d1, count6_d2, count6_d3 :  std_logic;
signal level6 :  std_logic_vector(89 downto 0);
signal count5, count5_d1, count5_d2, count5_d3 :  std_logic;
signal level5, level5_d1 :  std_logic_vector(89 downto 0);
signal count4, count4_d1, count4_d2 :  std_logic;
signal level4 :  std_logic_vector(88 downto 0);
signal count3, count3_d1, count3_d2 :  std_logic;
signal level3, level3_d1 :  std_logic_vector(80 downto 0);
signal count2, count2_d1 :  std_logic;
signal level2 :  std_logic_vector(76 downto 0);
signal count1, count1_d1 :  std_logic;
signal level1, level1_d1 :  std_logic_vector(74 downto 0);
signal count0 :  std_logic;
signal level0 :  std_logic_vector(73 downto 0);
signal sCount :  std_logic_vector(6 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            level7_d1 <=  level7;
            count6_d1 <=  count6;
            count6_d2 <=  count6_d1;
            count6_d3 <=  count6_d2;
            count5_d1 <=  count5;
            count5_d2 <=  count5_d1;
            count5_d3 <=  count5_d2;
            level5_d1 <=  level5;
            count4_d1 <=  count4;
            count4_d2 <=  count4_d1;
            count3_d1 <=  count3;
            count3_d2 <=  count3_d1;
            level3_d1 <=  level3;
            count2_d1 <=  count2;
            count1_d1 <=  count1;
            level1_d1 <=  level1;
         end if;
      end process;
   level7 <= I ;
   ----------------Synchro barrier, entering cycle 1----------------
   count6<= '1' when level7_d1(89 downto 26) = (89 downto 26=>'0') else '0';
   level6<= level7_d1(89 downto 0) when count6='0' else level7_d1(25 downto 0) & (63 downto 0 => '0');

   count5<= '1' when level6(89 downto 58) = (89 downto 58=>'0') else '0';
   level5<= level6(89 downto 0) when count5='0' else level6(57 downto 0) & (31 downto 0 => '0');

   ----------------Synchro barrier, entering cycle 2----------------
   count4<= '1' when level5_d1(89 downto 74) = (89 downto 74=>'0') else '0';
   level4<= level5_d1(89 downto 1) when count4='0' else level5_d1(73 downto 0) & (14 downto 0 => '0');

   count3<= '1' when level4(88 downto 81) = (88 downto 81=>'0') else '0';
   level3<= level4(88 downto 8) when count3='0' else level4(80 downto 0);

   ----------------Synchro barrier, entering cycle 3----------------
   count2<= '1' when level3_d1(80 downto 77) = (80 downto 77=>'0') else '0';
   level2<= level3_d1(80 downto 4) when count2='0' else level3_d1(76 downto 0);

   count1<= '1' when level2(76 downto 75) = (76 downto 75=>'0') else '0';
   level1<= level2(76 downto 2) when count1='0' else level2(74 downto 0);

   ----------------Synchro barrier, entering cycle 4----------------
   count0<= '1' when level1_d1(74 downto 74) = (74 downto 74=>'0') else '0';
   level0<= level1_d1(74 downto 1) when count0='0' else level1_d1(73 downto 0);

   O <= level0;
   sCount <= count6_d3 & count5_d3 & count4_d2 & count3_d2 & count2_d1 & count1_d1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                   RightShifter_28_by_max_27_F400_uid200
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter_28_by_max_27_F400_uid200 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(27 downto 0);
          S : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(54 downto 0)   );
end entity;

architecture arch of RightShifter_28_by_max_27_F400_uid200 is
signal level0 :  std_logic_vector(27 downto 0);
signal ps, ps_d1 :  std_logic_vector(4 downto 0);
signal level1 :  std_logic_vector(28 downto 0);
signal level2, level2_d1 :  std_logic_vector(30 downto 0);
signal level3 :  std_logic_vector(34 downto 0);
signal level4 :  std_logic_vector(42 downto 0);
signal level5 :  std_logic_vector(58 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level2_d1 <=  level2;
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   ----------------Synchro barrier, entering cycle 1----------------
   level3<=  (3 downto 0 => '0') & level2_d1 when ps_d1(2) = '1' else    level2_d1 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps_d1(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps_d1(4) = '1' else    level4 & (15 downto 0 => '0');
   R <= level5(58 downto 4);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_52_f400_uid204
--                    (IntAdderAlternative_52_F400_uid208)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_52_f400_uid204 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(51 downto 0);
          Y : in  std_logic_vector(51 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(51 downto 0)   );
end entity;

architecture arch of IntAdder_52_f400_uid204 is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(10 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(9 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(10 downto 0);
signal sum_l1_idx1 :  std_logic_vector(9 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(51 downto 42)) + ( "0" & Y(51 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
   sum_l0_idx1 <= s_sum_l0_idx1(9 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(10 downto 10);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(9 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(10 downto 10);
   R <= sum_l1_idx1(9 downto 0) & sum_l0_idx0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_62_f400_uid212
--                    (IntAdderAlternative_62_F400_uid216)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_62_f400_uid212 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(61 downto 0);
          Y : in  std_logic_vector(61 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(61 downto 0)   );
end entity;

architecture arch of IntAdder_62_f400_uid212 is
signal s_sum_l0_idx0 :  std_logic_vector(42 downto 0);
signal s_sum_l0_idx1, s_sum_l0_idx1_d1 :  std_logic_vector(20 downto 0);
signal sum_l0_idx0, sum_l0_idx0_d1 :  std_logic_vector(41 downto 0);
signal c_l0_idx0, c_l0_idx0_d1 :  std_logic_vector(0 downto 0);
signal sum_l0_idx1 :  std_logic_vector(19 downto 0);
signal c_l0_idx1 :  std_logic_vector(0 downto 0);
signal s_sum_l1_idx1 :  std_logic_vector(20 downto 0);
signal sum_l1_idx1 :  std_logic_vector(19 downto 0);
signal c_l1_idx1 :  std_logic_vector(0 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            s_sum_l0_idx1_d1 <=  s_sum_l0_idx1;
            sum_l0_idx0_d1 <=  sum_l0_idx0;
            c_l0_idx0_d1 <=  c_l0_idx0;
         end if;
      end process;
   --Alternative
   s_sum_l0_idx0 <= ( "0" & X(41 downto 0)) + ( "0" & Y(41 downto 0)) + Cin;
   s_sum_l0_idx1 <= ( "0" & X(61 downto 42)) + ( "0" & Y(61 downto 42));
   sum_l0_idx0 <= s_sum_l0_idx0(41 downto 0);
   c_l0_idx0 <= s_sum_l0_idx0(42 downto 42);
   sum_l0_idx1 <= s_sum_l0_idx1(19 downto 0);
   c_l0_idx1 <= s_sum_l0_idx1(20 downto 20);
   ----------------Synchro barrier, entering cycle 1----------------
   s_sum_l1_idx1 <=  s_sum_l0_idx1_d1 + c_l0_idx0_d1(0 downto 0);
   sum_l1_idx1 <= s_sum_l1_idx1(19 downto 0);
   c_l1_idx1 <= s_sum_l1_idx1(20 downto 20);
   R <= sum_l1_idx1(19 downto 0) & sum_l0_idx0_d1(41 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                          FPLog_16_46_0_F400_uid2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: F. de Dinechin, C. Klein  (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 21 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPLog_16_46_0_F400_uid2 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(16+46+2 downto 0);
          R : out  std_logic_vector(16+46+2 downto 0)   );
end entity;

architecture arch of FPLog_16_46_0_F400_uid2 is
   component LZOC_46_F400_uid4 is
      port ( clk, rst : in std_logic;
             I : in  std_logic_vector(45 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(5 downto 0)   );
   end component;

   component LeftShifter_24_by_max_24_F400_uid8 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component InvTable_0_10_11_F400_uid12 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(10 downto 0)   );
   end component;

   component IntAdder_59_f400_uid16 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(58 downto 0);
             Y : in  std_logic_vector(58 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(58 downto 0)   );
   end component;

   component IntAdder_59_f400_uid24 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(58 downto 0);
             Y : in  std_logic_vector(58 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(58 downto 0)   );
   end component;

   component IntAdder_50_f400_uid32 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(49 downto 0);
             Y : in  std_logic_vector(49 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(49 downto 0)   );
   end component;

   component IntAdder_50_f400_uid40 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(49 downto 0);
             Y : in  std_logic_vector(49 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(49 downto 0)   );
   end component;

   component IntSquarer_28_F400_uid48 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             R : out  std_logic_vector(55 downto 0)   );
   end component;

   component IntAdder_50_f400_uid52 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(49 downto 0);
             Y : in  std_logic_vector(49 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(49 downto 0)   );
   end component;

   component LogTable_0_10_74_F400_uid60 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(73 downto 0)   );
   end component;

   component LogTable_1_8_66_F400_uid76 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             Y : out  std_logic_vector(65 downto 0)   );
   end component;

   component IntAdder_74_f400_uid80 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(73 downto 0);
             Y : in  std_logic_vector(73 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(73 downto 0)   );
   end component;

   component LogTable_2_10_59_F400_uid88 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(58 downto 0)   );
   end component;

   component IntAdder_74_f400_uid92 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(73 downto 0);
             Y : in  std_logic_vector(73 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(73 downto 0)   );
   end component;

   component IntAdder_74_f400_uid100 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(73 downto 0);
             Y : in  std_logic_vector(73 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(73 downto 0)   );
   end component;

   component IntIntKCM_16_780414346020670_unsigned_F400_uid108 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(15 downto 0);
             R : out  std_logic_vector(65 downto 0)   );
   end component;

   component IntAdder_90_f400_uid188 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(89 downto 0);
             Y : in  std_logic_vector(89 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(89 downto 0)   );
   end component;

   component LZCShifter_90_to_74_counting_128_F400_uid196 is
      port ( clk, rst : in std_logic;
             I : in  std_logic_vector(89 downto 0);
             Count : out  std_logic_vector(6 downto 0);
             O : out  std_logic_vector(73 downto 0)   );
   end component;

   component RightShifter_28_by_max_27_F400_uid200 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(27 downto 0);
             S : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(54 downto 0)   );
   end component;

   component IntAdder_52_f400_uid204 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(51 downto 0);
             Y : in  std_logic_vector(51 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(51 downto 0)   );
   end component;

   component IntAdder_62_f400_uid212 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(61 downto 0);
             Y : in  std_logic_vector(61 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(61 downto 0)   );
   end component;

signal XExnSgn, XExnSgn_d1, XExnSgn_d2, XExnSgn_d3, XExnSgn_d4, XExnSgn_d5, XExnSgn_d6, XExnSgn_d7, XExnSgn_d8, XExnSgn_d9, XExnSgn_d10, XExnSgn_d11, XExnSgn_d12, XExnSgn_d13, XExnSgn_d14, XExnSgn_d15, XExnSgn_d16, XExnSgn_d17, XExnSgn_d18, XExnSgn_d19, XExnSgn_d20, XExnSgn_d21 :  std_logic_vector(2 downto 0);
signal FirstBit :  std_logic;
signal Y0, Y0_d1, Y0_d2 :  std_logic_vector(47 downto 0);
signal Y0h :  std_logic_vector(45 downto 0);
signal sR, sR_d1, sR_d2, sR_d3, sR_d4, sR_d5, sR_d6, sR_d7, sR_d8, sR_d9, sR_d10, sR_d11, sR_d12, sR_d13, sR_d14, sR_d15, sR_d16, sR_d17, sR_d18, sR_d19, sR_d20, sR_d21 :  std_logic;
signal absZ0, absZ0_d1, absZ0_d2, absZ0_d3, absZ0_d4 :  std_logic_vector(23 downto 0);
signal E, E_d1 :  std_logic_vector(15 downto 0);
signal absE, absE_d1, absE_d2, absE_d3, absE_d4, absE_d5, absE_d6, absE_d7, absE_d8, absE_d9, absE_d10 :  std_logic_vector(15 downto 0);
signal EeqZero, EeqZero_d1, EeqZero_d2, EeqZero_d3 :  std_logic;
signal lzo, lzo_d1, lzo_d2, lzo_d3, lzo_d4, lzo_d5, lzo_d6, lzo_d7, lzo_d8, lzo_d9, lzo_d10, lzo_d11, lzo_d12, lzo_d13, lzo_d14, lzo_d15, lzo_d16, lzo_d17 :  std_logic_vector(5 downto 0);
signal pfinal_s :  std_logic_vector(5 downto 0);
signal shiftval :  std_logic_vector(6 downto 0);
signal shiftvalinL :  std_logic_vector(4 downto 0);
signal shiftvalinR, shiftvalinR_d1, shiftvalinR_d2, shiftvalinR_d3, shiftvalinR_d4, shiftvalinR_d5, shiftvalinR_d6, shiftvalinR_d7, shiftvalinR_d8, shiftvalinR_d9, shiftvalinR_d10, shiftvalinR_d11, shiftvalinR_d12 :  std_logic_vector(4 downto 0);
signal doRR, doRR_d1, doRR_d2, doRR_d3 :  std_logic;
signal small, small_d1, small_d2, small_d3, small_d4, small_d5, small_d6, small_d7, small_d8, small_d9, small_d10, small_d11, small_d12, small_d13, small_d14, small_d15, small_d16, small_d17 :  std_logic;
signal small_absZ0_normd_full :  std_logic_vector(47 downto 0);
signal small_absZ0_normd, small_absZ0_normd_d1, small_absZ0_normd_d2, small_absZ0_normd_d3, small_absZ0_normd_d4, small_absZ0_normd_d5, small_absZ0_normd_d6, small_absZ0_normd_d7, small_absZ0_normd_d8, small_absZ0_normd_d9, small_absZ0_normd_d10, small_absZ0_normd_d11, small_absZ0_normd_d12 :  std_logic_vector(23 downto 0);
signal A0, A0_d1, A0_d2, A0_d3, A0_d4 :  std_logic_vector(9 downto 0);
signal InvA0 :  std_logic_vector(10 downto 0);
signal P0, P0_d1 :  std_logic_vector(58 downto 0);
signal Z1 :  std_logic_vector(48 downto 0);
signal A1, A1_d1, A1_d2 :  std_logic_vector(7 downto 0);
signal B1 :  std_logic_vector(40 downto 0);
signal ZM1, ZM1_d1 :  std_logic_vector(48 downto 0);
signal P1 :  std_logic_vector(56 downto 0);
signal Y1 :  std_logic_vector(57 downto 0);
signal EiY1 :  std_logic_vector(58 downto 0);
signal addXIter1 :  std_logic_vector(58 downto 0);
signal EiYPB1 :  std_logic_vector(58 downto 0);
signal Pp1 :  std_logic_vector(58 downto 0);
signal Z2 :  std_logic_vector(58 downto 0);
signal A2, A2_d1, A2_d2, A2_d3, A2_d4 :  std_logic_vector(9 downto 0);
signal B2 :  std_logic_vector(48 downto 0);
signal ZM2, ZM2_d1 :  std_logic_vector(43 downto 0);
signal P2 :  std_logic_vector(53 downto 0);
signal Y2 :  std_logic_vector(74 downto 0);
signal EiY2 :  std_logic_vector(49 downto 0);
signal addXIter2 :  std_logic_vector(49 downto 0);
signal EiYPB2 :  std_logic_vector(49 downto 0);
signal Pp2 :  std_logic_vector(49 downto 0);
signal Z3 :  std_logic_vector(49 downto 0);
signal Zfinal, Zfinal_d1, Zfinal_d2, Zfinal_d3, Zfinal_d4 :  std_logic_vector(49 downto 0);
signal squarerIn :  std_logic_vector(27 downto 0);
signal Z2o2_full :  std_logic_vector(55 downto 0);
signal Z2o2_full_dummy, Z2o2_full_dummy_d1, Z2o2_full_dummy_d2, Z2o2_full_dummy_d3, Z2o2_full_dummy_d4, Z2o2_full_dummy_d5 :  std_logic_vector(55 downto 0);
signal Z2o2_normal :  std_logic_vector(24 downto 0);
signal addFinalLog1pY :  std_logic_vector(49 downto 0);
signal Log1p_normal, Log1p_normal_d1 :  std_logic_vector(49 downto 0);
signal L0 :  std_logic_vector(73 downto 0);
signal S1, S1_d1, S1_d2 :  std_logic_vector(73 downto 0);
signal L1 :  std_logic_vector(65 downto 0);
signal sopX1, sopX1_d1, sopX1_d2 :  std_logic_vector(73 downto 0);
signal S2, S2_d1, S2_d2, S2_d3 :  std_logic_vector(73 downto 0);
signal L2 :  std_logic_vector(58 downto 0);
signal sopX2, sopX2_d1, sopX2_d2 :  std_logic_vector(73 downto 0);
signal S3, S3_d1 :  std_logic_vector(73 downto 0);
signal almostLog :  std_logic_vector(73 downto 0);
signal adderLogF_normalY :  std_logic_vector(73 downto 0);
signal LogF_normal :  std_logic_vector(73 downto 0);
signal absELog2 :  std_logic_vector(65 downto 0);
signal absELog2_pad :  std_logic_vector(89 downto 0);
signal LogF_normal_pad :  std_logic_vector(89 downto 0);
signal lnaddX :  std_logic_vector(89 downto 0);
signal lnaddY :  std_logic_vector(89 downto 0);
signal Log_normal :  std_logic_vector(89 downto 0);
signal E_normal :  std_logic_vector(6 downto 0);
signal Log_normal_normd, Log_normal_normd_d1 :  std_logic_vector(73 downto 0);
signal Z2o2_small_bs :  std_logic_vector(27 downto 0);
signal Z2o2_small_s :  std_logic_vector(54 downto 0);
signal Z2o2_small, Z2o2_small_d1 :  std_logic_vector(51 downto 0);
signal Z_small, Z_small_d1 :  std_logic_vector(51 downto 0);
signal Log_smallY :  std_logic_vector(51 downto 0);
signal nsRCin :  std_logic;
signal Log_small, Log_small_d1 :  std_logic_vector(51 downto 0);
signal E0_sub, E0_sub_d1 :  std_logic_vector(1 downto 0);
signal ufl, ufl_d1, ufl_d2 :  std_logic;
signal E_small :  std_logic_vector(15 downto 0);
signal Log_small_normd, Log_small_normd_d1 :  std_logic_vector(49 downto 0);
signal E0offset :  std_logic_vector(15 downto 0);
signal ER :  std_logic_vector(15 downto 0);
signal Log_g :  std_logic_vector(49 downto 0);
signal round :  std_logic;
signal fraX :  std_logic_vector(61 downto 0);
signal fraY :  std_logic_vector(61 downto 0);
signal EFR :  std_logic_vector(61 downto 0);
constant g: positive := 4;
constant log2wF: positive := 6;
constant pfinal: positive := 24;
constant sfinal: positive := 50;
constant targetprec: positive := 74;
constant wE: positive := 16;
constant wF: positive := 46;
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of InvTable_0_10_11_F400_uid12: component is "yes";
attribute rom_style of InvTable_0_10_11_F400_uid12: component is "block";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            XExnSgn_d1 <=  XExnSgn;
            XExnSgn_d2 <=  XExnSgn_d1;
            XExnSgn_d3 <=  XExnSgn_d2;
            XExnSgn_d4 <=  XExnSgn_d3;
            XExnSgn_d5 <=  XExnSgn_d4;
            XExnSgn_d6 <=  XExnSgn_d5;
            XExnSgn_d7 <=  XExnSgn_d6;
            XExnSgn_d8 <=  XExnSgn_d7;
            XExnSgn_d9 <=  XExnSgn_d8;
            XExnSgn_d10 <=  XExnSgn_d9;
            XExnSgn_d11 <=  XExnSgn_d10;
            XExnSgn_d12 <=  XExnSgn_d11;
            XExnSgn_d13 <=  XExnSgn_d12;
            XExnSgn_d14 <=  XExnSgn_d13;
            XExnSgn_d15 <=  XExnSgn_d14;
            XExnSgn_d16 <=  XExnSgn_d15;
            XExnSgn_d17 <=  XExnSgn_d16;
            XExnSgn_d18 <=  XExnSgn_d17;
            XExnSgn_d19 <=  XExnSgn_d18;
            XExnSgn_d20 <=  XExnSgn_d19;
            XExnSgn_d21 <=  XExnSgn_d20;
            Y0_d1 <=  Y0;
            Y0_d2 <=  Y0_d1;
            sR_d1 <=  sR;
            sR_d2 <=  sR_d1;
            sR_d3 <=  sR_d2;
            sR_d4 <=  sR_d3;
            sR_d5 <=  sR_d4;
            sR_d6 <=  sR_d5;
            sR_d7 <=  sR_d6;
            sR_d8 <=  sR_d7;
            sR_d9 <=  sR_d8;
            sR_d10 <=  sR_d9;
            sR_d11 <=  sR_d10;
            sR_d12 <=  sR_d11;
            sR_d13 <=  sR_d12;
            sR_d14 <=  sR_d13;
            sR_d15 <=  sR_d14;
            sR_d16 <=  sR_d15;
            sR_d17 <=  sR_d16;
            sR_d18 <=  sR_d17;
            sR_d19 <=  sR_d18;
            sR_d20 <=  sR_d19;
            sR_d21 <=  sR_d20;
            absZ0_d1 <=  absZ0;
            absZ0_d2 <=  absZ0_d1;
            absZ0_d3 <=  absZ0_d2;
            absZ0_d4 <=  absZ0_d3;
            E_d1 <=  E;
            absE_d1 <=  absE;
            absE_d2 <=  absE_d1;
            absE_d3 <=  absE_d2;
            absE_d4 <=  absE_d3;
            absE_d5 <=  absE_d4;
            absE_d6 <=  absE_d5;
            absE_d7 <=  absE_d6;
            absE_d8 <=  absE_d7;
            absE_d9 <=  absE_d8;
            absE_d10 <=  absE_d9;
            EeqZero_d1 <=  EeqZero;
            EeqZero_d2 <=  EeqZero_d1;
            EeqZero_d3 <=  EeqZero_d2;
            lzo_d1 <=  lzo;
            lzo_d2 <=  lzo_d1;
            lzo_d3 <=  lzo_d2;
            lzo_d4 <=  lzo_d3;
            lzo_d5 <=  lzo_d4;
            lzo_d6 <=  lzo_d5;
            lzo_d7 <=  lzo_d6;
            lzo_d8 <=  lzo_d7;
            lzo_d9 <=  lzo_d8;
            lzo_d10 <=  lzo_d9;
            lzo_d11 <=  lzo_d10;
            lzo_d12 <=  lzo_d11;
            lzo_d13 <=  lzo_d12;
            lzo_d14 <=  lzo_d13;
            lzo_d15 <=  lzo_d14;
            lzo_d16 <=  lzo_d15;
            lzo_d17 <=  lzo_d16;
            shiftvalinR_d1 <=  shiftvalinR;
            shiftvalinR_d2 <=  shiftvalinR_d1;
            shiftvalinR_d3 <=  shiftvalinR_d2;
            shiftvalinR_d4 <=  shiftvalinR_d3;
            shiftvalinR_d5 <=  shiftvalinR_d4;
            shiftvalinR_d6 <=  shiftvalinR_d5;
            shiftvalinR_d7 <=  shiftvalinR_d6;
            shiftvalinR_d8 <=  shiftvalinR_d7;
            shiftvalinR_d9 <=  shiftvalinR_d8;
            shiftvalinR_d10 <=  shiftvalinR_d9;
            shiftvalinR_d11 <=  shiftvalinR_d10;
            shiftvalinR_d12 <=  shiftvalinR_d11;
            doRR_d1 <=  doRR;
            doRR_d2 <=  doRR_d1;
            doRR_d3 <=  doRR_d2;
            small_d1 <=  small;
            small_d2 <=  small_d1;
            small_d3 <=  small_d2;
            small_d4 <=  small_d3;
            small_d5 <=  small_d4;
            small_d6 <=  small_d5;
            small_d7 <=  small_d6;
            small_d8 <=  small_d7;
            small_d9 <=  small_d8;
            small_d10 <=  small_d9;
            small_d11 <=  small_d10;
            small_d12 <=  small_d11;
            small_d13 <=  small_d12;
            small_d14 <=  small_d13;
            small_d15 <=  small_d14;
            small_d16 <=  small_d15;
            small_d17 <=  small_d16;
            small_absZ0_normd_d1 <=  small_absZ0_normd;
            small_absZ0_normd_d2 <=  small_absZ0_normd_d1;
            small_absZ0_normd_d3 <=  small_absZ0_normd_d2;
            small_absZ0_normd_d4 <=  small_absZ0_normd_d3;
            small_absZ0_normd_d5 <=  small_absZ0_normd_d4;
            small_absZ0_normd_d6 <=  small_absZ0_normd_d5;
            small_absZ0_normd_d7 <=  small_absZ0_normd_d6;
            small_absZ0_normd_d8 <=  small_absZ0_normd_d7;
            small_absZ0_normd_d9 <=  small_absZ0_normd_d8;
            small_absZ0_normd_d10 <=  small_absZ0_normd_d9;
            small_absZ0_normd_d11 <=  small_absZ0_normd_d10;
            small_absZ0_normd_d12 <=  small_absZ0_normd_d11;
            A0_d1 <=  A0;
            A0_d2 <=  A0_d1;
            A0_d3 <=  A0_d2;
            A0_d4 <=  A0_d3;
            P0_d1 <=  P0;
            A1_d1 <=  A1;
            A1_d2 <=  A1_d1;
            ZM1_d1 <=  ZM1;
            A2_d1 <=  A2;
            A2_d2 <=  A2_d1;
            A2_d3 <=  A2_d2;
            A2_d4 <=  A2_d3;
            ZM2_d1 <=  ZM2;
            Zfinal_d1 <=  Zfinal;
            Zfinal_d2 <=  Zfinal_d1;
            Zfinal_d3 <=  Zfinal_d2;
            Zfinal_d4 <=  Zfinal_d3;
            Z2o2_full_dummy_d1 <=  Z2o2_full_dummy;
            Z2o2_full_dummy_d2 <=  Z2o2_full_dummy_d1;
            Z2o2_full_dummy_d3 <=  Z2o2_full_dummy_d2;
            Z2o2_full_dummy_d4 <=  Z2o2_full_dummy_d3;
            Z2o2_full_dummy_d5 <=  Z2o2_full_dummy_d4;
            Log1p_normal_d1 <=  Log1p_normal;
            S1_d1 <=  S1;
            S1_d2 <=  S1_d1;
            sopX1_d1 <=  sopX1;
            sopX1_d2 <=  sopX1_d1;
            S2_d1 <=  S2;
            S2_d2 <=  S2_d1;
            S2_d3 <=  S2_d2;
            sopX2_d1 <=  sopX2;
            sopX2_d2 <=  sopX2_d1;
            S3_d1 <=  S3;
            Log_normal_normd_d1 <=  Log_normal_normd;
            Z2o2_small_d1 <=  Z2o2_small;
            Z_small_d1 <=  Z_small;
            Log_small_d1 <=  Log_small;
            E0_sub_d1 <=  E0_sub;
            ufl_d1 <=  ufl;
            ufl_d2 <=  ufl_d1;
            Log_small_normd_d1 <=  Log_small_normd;
         end if;
      end process;
   XExnSgn <=  X(wE+wF+2 downto wE+wF);
   FirstBit <=  X(wF-1);
   Y0 <= "1" & X(wF-1 downto 0) & "0" when FirstBit = '0' else "01" & X(wF-1 downto 0);
   Y0h <= Y0(wF downto 1);
   -- Sign of the result;
   sR <= '0'   when  (X(wE+wF-1 downto wF) = ('0' & (wE-2 downto 0 => '1')))  -- binade [1..2)
     else not X(wE+wF-1);                -- MSB of exponent
   absZ0 <=   Y0(wF-pfinal+1 downto 0)          when (sR='0') else
             ((wF-pfinal+1 downto 0 => '0') - Y0(wF-pfinal+1 downto 0));
   E <= (X(wE+wF-1 downto wF)) - ("0" & (wE-2 downto 1 => '1') & (not FirstBit));
   ----------------Synchro barrier, entering cycle 1----------------
   absE <= ((wE-1 downto 0 => '0') - E_d1)   when sR_d1 = '1' else E_d1;
   EeqZero <= '1' when E_d1=(wE-1 downto 0 => '0') else '0';
   ---------------- cycle 0----------------
   lzoc1: LZOC_46_F400_uid4  -- pipelineDepth=3 maxInDelay=6.38e-10
      port map ( clk  => clk,
                 rst  => rst,
                 I => Y0h,
                 O => lzo,
                 OZB => FirstBit);
   ---------------- cycle 3----------------
   ----------------Synchro barrier, entering cycle 4----------------
   pfinal_s <= "011000";
   shiftval <= ('0' & lzo_d1) - ('0' & pfinal_s); 
   shiftvalinL <= shiftval(4 downto 0);
   shiftvalinR <= shiftval(4 downto 0);
   doRR <= shiftval(log2wF); -- sign of the result
   small <= EeqZero_d3 and not(doRR);
   ---------------- cycle 4----------------
   -- The left shifter for the 'small' case
   small_lshift: LeftShifter_24_by_max_24_F400_uid8  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => small_absZ0_normd_full,
                 S => shiftvalinL,
                 X => absZ0_d4);
   ----------------Synchro barrier, entering cycle 5----------------
   small_absZ0_normd <= small_absZ0_normd_full(23 downto 0); -- get rid of leading zeroes
   ----------------Synchro barrier, entering cycle 0----------------
   ---------------- The range reduction box ---------------
   A0 <= X(45 downto 36);
   ----------------Synchro barrier, entering cycle 1----------------
   -- First inv table
   itO: InvTable_0_10_11_F400_uid12  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A0_d1,
                 Y => InvA0);
   ----------------Synchro barrier, entering cycle 2----------------
   P0 <= InvA0 * Y0_d2;

   ----------------Synchro barrier, entering cycle 3----------------
   Z1 <= P0_d1(48 downto 0);

   A1 <= Z1(48 downto 41);
   B1 <= Z1(40 downto 0);
   ZM1 <= Z1;
   ----------------Synchro barrier, entering cycle 4----------------
   P1 <= A1_d1*ZM1_d1;
   ----------------Synchro barrier, entering cycle 5----------------
    -- delay at multiplier output is 0
   ---------------- cycle 3----------------
   Y1 <= "1" & (7 downto 0 => '0') & Z1;
   EiY1 <= Y1 & (0 downto 0 => '0')  when A1(7) = '1'
     else  "0" & Y1;
   addXIter1 <= "0" & B1 & (16 downto 0 => '0');
   addIter1_1: IntAdder_59_f400_uid16  -- pipelineDepth=1 maxInDelay=8.6e-11
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0',
                 R => EiYPB1,
                 X => addXIter1,
                 Y => EiY1);

   ----------------Synchro barrier, entering cycle 4----------------
   Pp1 <= (0 downto 0 => '1') & not(P1 & (0 downto 0 => '0'));
   addIter2_1: IntAdder_59_f400_uid24  -- pipelineDepth=1 maxInDelay=1.059e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '1',
                 R => Z2,
                 X => EiYPB1,
                 Y => Pp1);

   ----------------Synchro barrier, entering cycle 5----------------
 -- the critical path at the adder output = 1.266e-09

   A2 <= Z2(58 downto 49);
   B2 <= Z2(48 downto 0);
   ZM2 <= Z2(58 downto 15);
   ----------------Synchro barrier, entering cycle 6----------------
   P2 <= A2_d1*ZM2_d1;
   ----------------Synchro barrier, entering cycle 7----------------
    -- delay at multiplier output is 0
   ---------------- cycle 5----------------
   Y2 <= "1" & (14 downto 0 => '0') & Z2;
   EiY2 <= (4 downto 0 => '0') & Y2(74 downto 30);
   addXIter2 <= "0" & B2;
   addIter1_2: IntAdder_50_f400_uid32  -- pipelineDepth=1 maxInDelay=1.266e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0',
                 R => EiYPB2,
                 X => addXIter2,
                 Y => EiY2);

   ----------------Synchro barrier, entering cycle 6----------------
   Pp2 <= (5 downto 0 => '1') & not(P2(53 downto 10));
   addIter2_2: IntAdder_50_f400_uid40  -- pipelineDepth=1 maxInDelay=1.266e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '1',
                 R => Z3,
                 X => EiYPB2,
                 Y => Pp2);

   ----------------Synchro barrier, entering cycle 7----------------
 -- the critical path at the adder output = 1.266e-09
   Zfinal <= Z3;
   --  Synchro between RR box and case almost 1
   squarerIn <= Zfinal(sfinal-1 downto sfinal-28) when doRR_d3='1'
                    else (small_absZ0_normd_d2 & (3 downto 0 => '0'));  
   squarer: IntSquarer_28_F400_uid48  -- pipelineDepth=4 maxInDelay=2.23272e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => Z2o2_full,
                 X => squarerIn);
   ----------------Synchro barrier, entering cycle 11----------------
   Z2o2_full_dummy <= Z2o2_full;
   Z2o2_normal <= Z2o2_full_dummy (55  downto 31);
   addFinalLog1pY <= (pfinal downto 0  => '1') & not(Z2o2_normal);
   addFinalLog1p_normalAdder: IntAdder_50_f400_uid52  -- pipelineDepth=1 maxInDelay=1.31672e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '1',
                 R => Log1p_normal,
                 X => Zfinal_d4,
                 Y => addFinalLog1pY);
   ----------------Synchro barrier, entering cycle 12----------------

   -- Now the log tables, as late as possible
   ----------------Synchro barrier, entering cycle 0----------------
   ----------------Synchro barrier, entering cycle 1----------------
   ----------------Synchro barrier, entering cycle 2----------------
   ----------------Synchro barrier, entering cycle 3----------------
   ----------------Synchro barrier, entering cycle 4----------------
   ----------------Synchro barrier, entering cycle 5----------------
   ----------------Synchro barrier, entering cycle 6----------------
   ----------------Synchro barrier, entering cycle 7----------------
   ----------------Synchro barrier, entering cycle 8----------------
   ----------------Synchro barrier, entering cycle 4----------------
   -- First log table
   ltO: LogTable_0_10_74_F400_uid60  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A0_d4,
                 Y => L0);
   ----------------Synchro barrier, entering cycle 5----------------
   S1 <= L0;
   lt1: LogTable_1_8_66_F400_uid76  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A1_d2,
                 Y => L1);
   sopX1 <= ((73 downto 66 => '0') & L1);
   ----------------Synchro barrier, entering cycle 6----------------
   ----------------Synchro barrier, entering cycle 7----------------
   adderS1: IntAdder_74_f400_uid80  -- pipelineDepth=1 maxInDelay=4.36e-10
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0' ,
                 R => S2,
                 X => S1_d2,
                 Y => sopX1_d2);

   ----------------Synchro barrier, entering cycle 8----------------
   ----------------Synchro barrier, entering cycle 9----------------
   lt2: LogTable_2_10_59_F400_uid88  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => A2_d4,
                 Y => L2);
   sopX2 <= ((73 downto 59 => '0') & L2);
   ----------------Synchro barrier, entering cycle 10----------------
   ----------------Synchro barrier, entering cycle 11----------------
   adderS2: IntAdder_74_f400_uid92  -- pipelineDepth=1 maxInDelay=4.36e-10
      port map ( clk  => clk,
                 rst  => rst,
                 Cin =>  '0' ,
                 R => S3,
                 X => S2_d3,
                 Y => sopX2_d2);

   ----------------Synchro barrier, entering cycle 12----------------
   ----------------Synchro barrier, entering cycle 13----------------
   almostLog <= S3_d1;
   adderLogF_normalY <= ((targetprec-1 downto sfinal => '0') & Log1p_normal_d1);
   adderLogF_normal: IntAdder_74_f400_uid100  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => '0',
                 R => LogF_normal,
                 X => almostLog,
                 Y => adderLogF_normalY);
   ----------------Synchro barrier, entering cycle 14----------------
   ----------------Synchro barrier, entering cycle 11----------------
   Log2KCM: IntIntKCM_16_780414346020670_unsigned_F400_uid108  -- pipelineDepth=3 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => absELog2,
                 X => absE_d10);
   ----------------Synchro barrier, entering cycle 14----------------
   absELog2_pad <=   absELog2 & (targetprec-wF-g-1 downto 0 => '0');       
   LogF_normal_pad <= (wE-1  downto 0 => LogF_normal(targetprec-1))  & LogF_normal;
   lnaddX <= absELog2_pad;
   lnaddY <= LogF_normal_pad when sR_d14='0' else not(LogF_normal_pad); 
   lnadder: IntAdder_90_f400_uid188  -- pipelineDepth=2 maxInDelay=1.49e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => sR_d14,
                 R => Log_normal,
                 X => lnaddX,
                 Y => lnaddY);

   ----------------Synchro barrier, entering cycle 16----------------
   final_norm: LZCShifter_90_to_74_counting_128_F400_uid196  -- pipelineDepth=4 maxInDelay=1.89472e-09
      port map ( clk  => clk,
                 rst  => rst,
                 Count => E_normal,
                 I => Log_normal,
                 O => Log_normal_normd);
   Z2o2_small_bs <= Z2o2_full_dummy_d5(55 downto 28);
   ao_rshift: RightShifter_28_by_max_27_F400_uid200  -- pipelineDepth=1 maxInDelay=5.3072e-10
      port map ( clk  => clk,
                 rst  => rst,
                 R => Z2o2_small_s,
                 S => shiftvalinR_d12,
                 X => Z2o2_small_bs);
   ---------------- cycle 17----------------
   -- output delay at shifter output is 1.93344e-09
     -- send the MSB to position pfinal
   Z2o2_small <=  (pfinal-1 downto 0  => '0') & Z2o2_small_s(54 downto 27);
   -- mantissa will be either Y0-z^2/2  or  -Y0+z^2/2,  depending on sR  
   Z_small <= small_absZ0_normd_d12 & (27 downto 0 => '0');
   ----------------Synchro barrier, entering cycle 18----------------
   Log_smallY <= Z2o2_small_d1 when sR_d18='1' else not(Z2o2_small_d1);
   nsRCin <= not ( sR_d18 );
   log_small_adder: IntAdder_52_f400_uid204  -- pipelineDepth=1 maxInDelay=4.4472e-10
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => nsRCin,
                 R => Log_small,
                 X => Z_small_d1,
                 Y => Log_smallY);

   ----------------Synchro barrier, entering cycle 19----------------
 -- critical path here is 8.98e-10
   -- Possibly subtract 1 or 2 to the exponent, depending on the LZC of Log_small
   E0_sub <=   "11" when Log_small(wF+g+1) = '1'
          else "10" when Log_small(wF+g+1 downto wF+g) = "01"
          else "01" ;
   -- The smallest log will be log(1+2^{-wF}) \approx 2^{-wF}  = 2^-46
   -- The smallest representable number is 2^{1-2^(wE-1)} = 2^-32767
   -- No underflow possible
   ufl <= '0';
   ----------------Synchro barrier, entering cycle 20----------------
   E_small <=  ("0" & (wE-2 downto 2 => '1') & E0_sub_d1)  -  ((wE-1 downto 6 => '0') & lzo_d17) ;
   Log_small_normd <= Log_small_d1(wF+g+1 downto 2) when Log_small_d1(wF+g+1)='1'
           else Log_small_d1(wF+g downto 1)  when Log_small_d1(wF+g)='1'  -- remove the first zero
           else Log_small_d1(wF+g-1 downto 0)  ; -- remove two zeroes (extremely rare, 001000000 only)
   E0offset <= "1000000000001110"; -- E0 + wE 
   ER <= E_small(15 downto 0) when small_d16='1'
      else E0offset - ((15 downto 7 => '0') & E_normal);
   ---------------- cycle 20----------------
   Log_g <=  Log_small_normd(wF+g-2 downto 0) & "0" when small_d16='1'           -- remove implicit 1
      else Log_normal_normd(targetprec-2 downto targetprec-wF-g-1 );  -- remove implicit 1
   round <= Log_g(g-1) ; -- sticky is always 1 for a transcendental function 
   -- if round leads to a change of binade, the carry propagation magically updates both mantissa and exponent
   fraX <= (ER & Log_g(wF+g-1 downto g)) ; 
   fraY <= ((wE+wF-1 downto 1 => '0') & round); 
   finalRoundAdder: IntAdder_62_f400_uid212  -- pipelineDepth=1 maxInDelay=6.1672e-10
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => '0',
                 R => EFR,
                 X => fraX,
                 Y => fraY);
   ----------------Synchro barrier, entering cycle 21----------------
   R(wE+wF+2 downto wE+wF) <= "110" when ((XExnSgn_d21(2) and (XExnSgn_d21(1) or XExnSgn_d21(0))) or (XExnSgn_d21(1) and XExnSgn_d21(0))) = '1' else
                              "101" when XExnSgn_d21(2 downto 1) = "00"  else
                              "100" when XExnSgn_d21(2 downto 1) = "10"  else
                              "00" & sR_d21 when (((Log_normal_normd_d1(targetprec-1)='0') and (small_d17='0')) or ( (Log_small_normd_d1 (wF+g-1)='0') and (small_d17='1'))) or (ufl_d2 = '1') else
                               "01" & sR_d21;
   R(wE+wF-1 downto 0) <=  EFR;
end architecture;

--------------------------------------------------------------------------------
--               TestBench_FPLog_16_46_0_F400_uid2_F400_uid220
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Cristian Klein, Nicolas Brunie (2007-2010)
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity TestBench_FPLog_16_46_0_F400_uid2_F400_uid220 is
end entity;

architecture behavorial of TestBench_FPLog_16_46_0_F400_uid2_F400_uid220 is
   component FPLog_16_46_0_F400_uid2 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(16+46+2 downto 0);
             R : out  std_logic_vector(16+46+2 downto 0)   );
   end component;
   signal X :  std_logic_vector(64 downto 0);
   signal R :  std_logic_vector(16+46+2 downto 0);
   signal clk :  std_logic;
   signal rst :  std_logic;

   -- FP compare function (found vs. real)
   function fp_equal(a : std_logic_vector; b : std_logic_vector) return boolean is
   begin
      if b(b'high downto b'high-1) = "01" then
         return a = b;
      elsif b(b'high downto b'high-1) = "11" then
         return (a(a'high downto a'high-1)=b(b'high downto b'high-1));
      else
         return a(a'high downto a'high-2) = b(b'high downto b'high-2);
      end if;
   end;



 -- converts std_logic into a character
   function chr(sl: std_logic) return character is
      variable c: character;
   begin
      case sl is
         when 'U' => c:= 'U';
         when 'X' => c:= 'X';
         when '0' => c:= '0';
         when '1' => c:= '1';
         when 'Z' => c:= 'Z';
         when 'W' => c:= 'W';
         when 'L' => c:= 'L';
         when 'H' => c:= 'H';
         when '-' => c:= '-';
      end case;
      return c;
   end chr;
   -- converts bit to std_logic (1 to 1)
   function to_stdlogic(b : bit) return std_logic is
       variable sl : std_logic;
   begin
      case b is 
         when '0' => sl := '0';
         when '1' => sl := '1';
      end case;
      return sl;
   end to_stdlogic;
   -- converts std_logic into a string (1 to 1)
   function str(sl: std_logic) return string is
    variable s: string(1 to 1);
    begin
      s(1) := chr(sl);
      return s;
   end str;
   -- converts std_logic_vector into a string (binary base)
   -- (this also takes care of the fact that the range of
   --  a string is natural while a std_logic_vector may
   --  have an integer range)
   function str(slv: std_logic_vector) return string is
      variable result : string (1 to slv'length);
      variable r : integer;
   begin
      r := 1;
      for i in slv'range loop
         result(r) := chr(slv(i));
         r := r + 1;
      end loop;
      return result;
   end str;




   -- test isZero
   function iszero(a : std_logic_vector) return boolean is
   begin
      return  a = (a'high downto 0 => '0');
   end;


   -- FP IEEE compare function (found vs. real)
   function fp_equal_ieee(a : std_logic_vector; b : std_logic_vector; we : integer; wf : integer) return boolean is
   begin
      if a(wf+we downto wf) = b(wf+we downto wf) and b(we+wf-1 downto wf) = (we downto 1 => '1') then
         if iszero(b(wf-1 downto 0)) then return  iszero(a(wf-1 downto 0));
         else return not iszero(a(wf - 1 downto 0));
         end if;
      else
         return a(a'high downto 0) = b(b'high downto 0);
      end if;
   end;

   -- FP subtypes for casting
   subtype fp65 is std_logic_vector(64 downto 0);
begin
   test: FPLog_16_46_0_F400_uid2  -- pipelineDepth=21 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => R,
                 X => X);
   -- Ticking clock signal
   process
   begin
      clk <= '0';
      wait for 5 ns;
      clk <= '1';
      wait for 5 ns;
   end process;

   -- Reading the input from a file 
   process
      variable inline : line; 
      variable counter : integer := 1;
      variable errorCounter : integer := 0;
      variable possibilityNumber : integer := 0;
      variable localErrorCounter : integer := 0;
      variable tmpChar : character;
      file inputsFile : text is "test.input"; 
      variable V_X : bit_vector(64 downto 0);
      variable V_R : bit_vector(64 downto 0);
   begin
      -- Send reset
      rst <= '1';
      wait for 10 ns;
      rst <= '0';
      while not endfile(inputsFile) loop
          -- positionning inputs
         readline(inputsFile,inline);
         read(inline ,V_X);
         read(inline,tmpChar);
         X <= to_stdlogicvector(V_X);
         readline(inputsFile,inline);
         wait for 10 ns;
      end loop;
      wait for 10000 ns; -- wait for simulation to finish
   end process;
          -- verifying the corresponding output
         process
      variable inline0 : line; 
      variable inline : line; 
      variable counter : integer := 1;
      variable errorCounter : integer := 0;
      variable possibilityNumber : integer := 0;
      variable localErrorCounter : integer := 0;
      variable tmpChar : character;
      file inputsFile : text is "test.input"; 
      variable V_R : bit_vector(64 downto 0);
      variable expected_R: string (1 to 1000);
      variable expected_size_R : integer;
   begin
          wait for 10 ns;
      wait for 210 ns; -- wait for pipeline to flush
      while not endfile(inputsFile) loop
          -- positionning inputs
         readline(inputsFile,inline0);
         readline(inputsFile,inline);
         read(inline, possibilityNumber);
         localErrorCounter := 0; -- 0 means error
         read(inline,tmpChar);
         expected_size_R := inline'Length;
         expected_R := inline.all & (expected_size_R+1 to 1000 => ' ');
         if possibilityNumber = 0 then
            localErrorCounter := 0;
         elsif possibilityNumber = 1 then 
            read(inline ,V_R);
            if not fp_equal(fp65'(R) ,to_stdlogicvector(V_R)) then 
               assert false report("Line " & integer'image(counter) & " of input file, incorrect output for R: " & lf & "  expected value: " & expected_R(1 to expected_size_R) & lf & "          result: " & str(R)) ;
               errorCounter := errorCounter + 1; -- incrementing global error counter
            end if;
         else
            for i in possibilityNumber downto 1 loop 
               read(inline ,V_R);
               read(inline,tmpChar);
               if fp_equal(fp65'(R) ,to_stdlogicvector(V_R))   then localErrorCounter := 1; end if; 
            end loop;
             if (localErrorCounter = 0) then 
               errorCounter := errorCounter + 1; -- incrementing global error counter
               assert false report("Line " & integer'image(counter) & " of input file, incorrect output for R: " & lf & " expected values: " & expected_R(1 to expected_size_R) & lf & "          result: " & str(R)) ;
            end if;
         end if;
          wait for 10 ns; -- wait for pipeline to flush
         counter := counter + 2;
      end loop;
      report (integer'image(errorCounter) & " error(s) encoutered.");
      report "End of simulation" severity note;
   end process;

end architecture;

