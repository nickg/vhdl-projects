-- *********************************************************************/ 
-- Copyright 2006 Actel Corporation.  All rights reserved.
-- IP Solutions Group
--  
-- File:  EDAC NETLIST
--     
-- Description: EDAC
--                
--
-- Rev: 1.0  01Jul02 HC  : Initial Code  
-- Rev: 1.3  17May06 IPB : Fixed Simultanous read/write SARS
-- Rev: 1.4  01Jun06 IPB : Removed W2R port
-- Rev: 1.5  06Jun06 IPB : fixed SLOWDOWN issue SAR	56406
--
-- Notes:
--
--
-- *********************************************************************/ 
--
--
--
library IEEE,axcelerator;

use IEEE.std_logic_1164.all;
use axcelerator.components.all;

package CONV_PACK_edaci is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_edaci;

library IEEE,axcelerator;

use IEEE.std_logic_1164.all;
use axcelerator.components.all;

use work.CONV_PACK_edaci.all;

entity edaci is

   port( waddr, raddr, wdata : in std_logic_vector (11 downto 0);  rdata : out 
         std_logic_vector (11 downto 0);  tmout : in std_logic_vector (41 
         downto 0);  rds : in std_logic_vector (3 downto 0);  wp : in 
         std_logic_vector (5 downto 0);  rp : out std_logic_vector (5 downto 0)
         ;  caddr, axwaddr, axraddr : out std_logic_vector (11 downto 0);  
         axwdata : out std_logic_vector (17 downto 0);  axrdata : in 
         std_logic_vector (17 downto 0);  clk, we, re, rstn, stop_scrub, bypass
         : in std_logic;  slowdown, scrub_corrected, error, scrub_done, 
         tmoutflg, correctable, axwe, axre : out std_logic);

end edaci;

architecture SYN_DEF_ARCH of edaci is

signal VXXXXXXXX, XXXDXXXXXXXXXXXXXXXX, XXDDXXXXXQ, XXXXXXXXXXXXXXXXX, 
   XXDXXXXXX, XXDDXXXXXJ, XXXDXXXXDXXXXYXXXXX, 
   XXXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXX, XXYPXXXXXX, XXDDXXXXXL, XXDDXXXXX, 
   XXXXXXDXXXX, XXDDXXXXXW, XXDDXXXXXXF, XXXXXXXXXXXXXXXXXF, XXDDXXXXXX, 
   XXDDXXXXXF, XXDDXXXXXV, XXDDXXXXXK, XXDDXXXXXH, XXDDXXXXXP, XXDXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXL, XXDXXXXXXXXXXF, XXDXXXXXXXXXXH, XXDXXXXXXXXXXXXXXP, 
   XXDXXXXXXXXXXJ, XXDXXXXXXXX, XXDXXXXXXXXXXK, XXDXXXXXXXXXXL, XXDXXXXXXXXXXP,
   XXDXXXXXXXXXXQ, XXDXXXXXXXXXXV, XXDXXXXXXXXXXW, XXDXXXXXXXXXXXXXXQ, 
   XXDXXXXXXXXF, XXDXXXXXXXXXXFD, XXDXXXXXXXXXXXXXXV, XXDXXXXXXXXXXFF, 
   XXDXXXXXXXXXXFH, XXDXXXXXXXXXXFJ, XXDXXXXXXXXXXFK, XXDXXXXXXXXXXFL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXFP, XXDXXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXFQ, XXDXXXXXXXXXXFV, XXDXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXFW, 
   XXDXXXXXXXXXXHD, XXDXXXXXXXXXXHF, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXDXDXXXXXXXXV, XXDXXXXXXXXXXXDXDXXXXXXH, 
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXDXD, 
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXX, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXDXXXXXYXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXXXX, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXDXXXXXYXXXXXXXXXXXXXF, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, XXDXXXXDXXXXXYXXXXXXXXXXXXXH, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, XXDXXXXDXXXXXXXXXXXXLXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXFD, XXDXXXXDXXXXXYXXXXXH, XXDXXXXDXXXXXYXXXXXJ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, XXDXXXXDXXXXXYXXXXXXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXF, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, XXDXXXXDXXXXXYXXXXXXXXXXXXXJ, 
   XXDXXXXDXXXXXXXXXX, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, 
   XXDXXXXDXXXXXXXX, XXDXXXXDXXXXXXXXF, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, XXDXXXXDXXXXXYXXXXXK, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXF,
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, XXDXXXXDXXXXXYXXXXXL, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXK, XXDXXXXDXXXXXXXXH, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXL, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXP, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXFP, XXDXXXXXXXXXXYXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXLXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXH, XXDXXXXXXXXXXXXXXFF, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXDDXXLXXXXXXX, XXDXXXXXXXXXXY, 
   XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, XXDXXXXXXXXXXXXXXDDXXLXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXFQ, XXDXXXXXXXXXXYXXX, XXDXXXXXXXXXXXXXXXFV, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXF, 
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, XXDXXXXXXXXXXYXXF, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXJ, XXDXXXXXXXXXXXXXXXXXXXXLXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXDDXXLXXXXXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, XXDXXXXXXXXXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXF
   , XXDXXXXXXXXXXXXXXXXXXXXXXQXXXX, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXJ, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXDDXLDXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXF, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXK, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXFF, XXDXXXXXXXXXXXXXXXFW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXHD, 
   XXDXXXXXXXXXXXXXXFH, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, XXDXXXXXXXXXXXXXXFJ
   , XXDXXXXXXXXXXYXXH, XXDXXXXXXXXXXXFXXXXLXXDX, XXDXXXXXXXXXXXXXXXXXXXXQ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJJ, XXDXXXXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXDDXXXXXFD, XXDXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXDDXXLXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXJK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXH, XXDXXXXXXXXXXXXXXFK, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXXXXXDDXXXXXFF, 
   XXDXXXXXXXXXXXXXXXHF, XXDXXXXXXXXXXXXXXXHH, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXJ,
   XXDXXXXXXXXXXXXXXXDDXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXK, XXDXXXXXXXXXXXXXXXXXXXXLXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXV, XXDXXXXXXXXXXXXXXDDXXLXXXXXXXX, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXK, XXDXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXP, XXDXXXXXXXXXXXXXXXXXXXXLXXXQ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, 
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXFL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, XXDXXXXXXXXXXXXXXDDXXLXXF, 
   XXDXXXXXXXXXXXXXXXHJ, XXDXXXXXXXXXXXXXXDDXXLXXXXXXXXF, XXDXXXXXXXXXXXXXXXHK,
   XXDXXXXXXXXXXYXXJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXQ, XXDXXXXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXDDXXXXXFH, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXW, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFD, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, 
   XXDXXXXXXXXXXXXXXXHL, XXDXXXXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXXXLXXXFF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXV, XXDXXXXXXXXXXXXWXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFH, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXW, 
   XXDXXXXXXXXXXXXXXDDXXLXXXXXXXJ, XXDXXXXXXXXXXXXXXXHP, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, XXDXXXXXXXXXXYXXK, 
   XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXHQ, 
   XXDXXXXXXXXXXXXXXDDXXLXXH, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFD, 
   XXDXXXXXXXXXXXXXXDDXXLXXJ, XXDXXXXXXXXXXXXXXDDXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXDDXXXXXFJ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXLXXXFJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFK, XXDXXXXXXXXXXXXXXXWXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXXXXXXWXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXFLXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, 
   XXDXXXXXXXXXXXXXXXHV, XXDXXXXXXXXXXYXXL, XXDXXXXXXXXXXXXXXDDXXLXXX, 
   XXDXXXXXXXXXXXXXXDDXXLXXK, XXDXXXXXXXXXXYXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, XXDXXXXXXXXXXXXXXXXXXXXLXXXFL, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFP, XXDXXXXXXXXXXXXXXDDXXLXXL, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFQ, XXDXXXXXXXXXXXXXXDDXXLXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH, 
   XXDXXXXXXXXXXXXXXDDXLDXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXF, 
   XXDXXXXXXXXXXYXXP, XXDXXXXXXXXXXXXXXDDXXXXXFK, XXDXXXXXXXXXXXXXXXHW, 
   XXDXXXXXXXXXXXXXXDDXXLXXXF, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFV, XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXJD, XXDXXXXXXXXXXXXXXXXXXXXLXXXFW, XXDXXXXXXXXXXXXXXXFLXX,
   XXDXXXXXXXXXXXXXXXXXP, XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXYXXXH, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXP, XXDXXXXXXXXXXXXXXXXXXXXLXXXHD, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXL, XXDXXXXXXXXXXXXXXXXXXXXLXXXHF, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHH, XXDXXXXXXXXXXXXXXXXXQ, 
   XXDXXXXXXXXXXXXXXDDXXLXXQ, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXQ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFH, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXP, XXDXXXXXXXXXXXXXXXXXXXXLXXXHJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXJF, 
   XXDXXXXXXXXXXXXXXFP, XXDXXXXXXXXXXXXXXDDXXLXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHK, XXDXXXXXXXXXXXXXXDDXXLXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXHL, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFK, XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXJL, 
   XXDXXXXXXXXXXXXXXDDXXLXXW, XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHP, XXDXXXXXXXXXXXXXXXXXXXXLXXXHQ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXHV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, XXDXXXXXXXXXXXXXXXXXXXXLXXXHW, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFL, XXDXXXXXXXXXXXXXXXJH, 
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, XXDXXXXXXXXXXYXXQ, XXDXXXXXXXXXXXXXXDDXXXXXFL
   , XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXQ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, 
   XXDXXXXXXXXXXXXXXDDXXLXXXXXXXL, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFP, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXJD, XXDXXXXXXXXXXXXXXXXXXXXLXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF
   , XXDXXXXXXXXXXXXXXXXXV, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXXXXXXJJ, 
   XXDXXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFQ, 
   XXDXXXXXXXXXXXXXXDDXXLXXXXXXXP, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFV, 
   XXDXXXXXXXXXXXXXXXJK, XXDXXXXXXXXXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFW, 
   XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHD, 
   XXDXXXXXXXXXXXXXXDDXXLXXXXXXXQ, XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXDDXXF, XXDXXXXXXXXXXXXXXXJL, XXDXXXXXXXXXXYXXV, 
   XXDXXXXXXXXXXXXXXFQ, XXDXXXXXXXXXXXXXXXXXXXXLXXP, XXDXXXXXXXXXXXXXXXJP, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, XXDXXXXXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXXXXXXXXXXXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXQ, XXDXXXXXXXXXXXXXXXXXXXXLXXXJF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHH, XXDXXXXXXXXXXXXXXXJQ, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXV, XXDXXXXXXXXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXV, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXQ, XXDXXXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJP, XXDXXXXXXXXXXYXXW, XXDXXXXXXXXXXXXXXFV, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHJ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, 
   XXDXXXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXFF, XXDXXXXXXXXXXXXXXXXXXXXLXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHK, XXDXXXXXXXXXXXXXXDDXXX, 
   XXDXXXXXXXXXXXXXXXJV, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, 
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXQ, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXW, XXDXXXXXXXXXXXXXXFW, 
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXW, XXDXXXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXW, XXDXXXXXXXXXXYXXXJ : std_logic;

begin
   caddr <= ( XXDDXXXXXX, XXDDXXXXXXF, XXDDXXXXX, XXDDXXXXXF, XXDDXXXXXH, 
      XXDDXXXXXJ, XXDDXXXXXK, XXDDXXXXXL, XXDDXXXXXP, XXDDXXXXXQ, XXDDXXXXXV, 
      XXDDXXXXXW );
   scrub_done <= XXXXXXDXXXX;
   
   XVXXX : VCC port map( Y => VXXXXXXXX);
   XXXXXXXXXXXXXXX : CM8INV port map( A => XXXDXXXXXXXXXXXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXX);
   XXXXXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => VXXXXXXXX, D2 => 
                           XXXXXXXXXXXXXXXXXF, D3 => XXDXXXXXX, S00 => 
                           XXXXXXXXXXXXXXXXXF, S01 => 
                           XXXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXX, S10 => 
                           XXXDXXXXDXXXXYXXXXX, S11 => XXDXXXXXX, Y => 
                           correctable);
   XXXDX : GND port map( Y => XXDXXXXXX);
   XYPXXXXX : BUFF port map( A => bypass, Y => XXYPXXXXXX);
   XXXXXXXXXXF : CM8 port map( D0 => XXXXXXXXXXXXXXXXX, D1 => XXDXXXXXX, D2 => 
                           XXDXXXXXX, D3 => VXXXXXXXX, S00 => XXXXXXXXXXXXXXXXX
                           , S01 => XXXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXX, S10 => 
                           XXXDXXXXDXXXXYXXXXX, S11 => XXDXXXXXX, Y => error);
   XXXXXXXXXXXXXXXF : CM8INV port map( A => XXXDXXXXXXXXXXXXXXXX, Y => 
                           XXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXDXDXXXXXXXX : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXV, C => wdata(0), D => 
                           wdata(3), Y => XXDXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXDXDXXXXXXXXF : CM8 port map( D0 => wdata(9), D1 => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXX, D3 => wdata(9)
                           , S00 => wdata(1), S01 => VXXXXXXXX, S10 => wdata(3)
                           , S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXDXDXXXXXXXXH : XOR2 port map( A => wdata(10), B => wdata(8), Y
                           => XXDXXXXXXXXXXXDXDXXXXXXXXV);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXX : CM8INV port map( A => wdata(9), Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXDXDXX : XOR4 port map( A => wdata(4), B => wdata(6), C => 
                           wdata(0), D => wdata(2), Y => XXDXXXXXXXXXXXXXXXDXD)
                           ;
   XXDXXXXXXXXXXXDXDXXXXXX : XOR2 port map( A => XXDXXXXXXXXXXXXXXXDXD, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXV, Y => XXDXXXXXXXXXXXXXXW)
                           ;
   XXDXXXXXXXXXXXDXDXXXXXXXXJ : XOR2 port map( A => wdata(11), B => 
                           XXDXXXXXXXXXXXDXDXXXXXXH, Y => XXDXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXDXDXXXXXXXXK : XOR2 port map( A => wdata(7), B => wdata(5), Y 
                           => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXDXDXXXXXXXXL : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX, B => wdata(1), C =>
                           wdata(2), D => wdata(8), Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXH);
   XXDXXXXXXXXXXXDXDXXXXXXXXP : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF, B => wdata(5), C 
                           => wdata(6), D => wdata(11), Y => XXDXXXXXXXXXXXXXXQ
                           );
   XXDXXXXXXXXXXXDXDXXXXXXF : CM8 port map( D0 => wdata(11), D1 => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXX, D3 => wdata(11),
                           S00 => XXDXXXXXXXXXXXXXXXDXD, S01 => VXXXXXXXX, S10 
                           => wdata(9), S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXDXDXXXXXXXXQ : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF, B => wdata(4), C 
                           => wdata(7), D => wdata(10), Y => XXDXXXXXXXXXXXXXXV
                           );
   XXDXXXXXXXXXXXDXDXXXXXXXXXXX : CM8INV port map( A => wdata(11), Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXDXXXXXXXXXX, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => axrdata(17), Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXK, D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, D2 => 
                           XXDXXXXXX, D3 => VXXXXXXXX, S00 => axrdata(1), S01 
                           => VXXXXXXXX, S10 => XXDXXXXDXXXXXXXXF, S11 => 
                           XXDXXXXXXXX, Y => XXDXXXXXXXXXXFH);
   XXDXXXXDXXXXXYXXXXXXX : XOR4 port map( A => axrdata(16), B => axrdata(13), C
                           => axrdata(15), D => XXDXXXXDXXXXXYXXXXXXXXXXXXXH, Y
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXYXXXXXXXF : XOR4 port map( A => axrdata(12), B => axrdata(11), 
                           C => axrdata(5), D => XXDXXXXDXXXXXYXXXXXXXXXXXXXH, 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXP);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => XXDXXXXXXXXXXK, Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => XXDXXXXXXXXF, Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXDXXXXXXXXXX, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => XXDXXXXXXXXXXK, Y
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXDXXXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, S00 => 
                           XXDXXXXXXXXXXF, S01 => XXDXXXXXXXXXXK, S10 => 
                           axrdata(12), S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXFP)
                           ;
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => axrdata(9), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D2 => 
                           axrdata(9), D3 => axrdata(9), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXXXXXXXFL, S10 =>
                           XXDXXXXDXXXXXYXXXXXH, S11 => XXDXXXXDXXXXXXXXH, Y =>
                           XXDXXXXXXXXXXW);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXH : AND2A port map( A => 
                           XXDXXXXDXXXXXYXXXXXL, B => XXDXXXXDXXXXXYXXXXXK, Y 
                           => XXDXXXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXJ, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S00 => 
                           XXDXXXXXXXXXXK, S01 => XXDXXXXXXXXXXFL, S10 => 
                           axrdata(4), S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXHD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXJ : AND2A port map( A => 
                           XXDXXXXDXXXXXYXXXXXK, B => XXDXXXXDXXXXXYXXXXXL, Y 
                           => XXDXXXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXF, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, S00 => 
                           XXDXXXXXXXXXXK, S01 => XXDXXXXXXXXXXFL, S10 => 
                           axrdata(5), S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D2 => 
                           VXXXXXXXX, D3 => XXDXXXXXXXXF, S00 => XXDXXXXXXXXXXJ
                           , S01 => XXDXXXXXXXXXXFL, S10 => axrdata(13), S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXFK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXK, D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXXX, D3 => VXXXXXXXX, S00 => axrdata(0), S01 
                           => VXXXXXXXX, S10 => XXDXXXXDXXXXXXXX, S11 => 
                           XXDXXXXXXXX, Y => XXDXXXXXXXXXXP);
   XXDXXXXDXXXXXYXXXXXXXXX : XOR4 port map( A => axrdata(10), B => axrdata(12),
                           C => axrdata(6), D => axrdata(8), Y => 
                           XXDXXXXDXXXXXYXXXXXXXFD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXL : CM8 port map( D0 => axrdata(8), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D2 => 
                           axrdata(8), D3 => axrdata(8), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXDXXXXXXXXXX, S10
                           => XXDXXXXDXXXXXYXXXXXJ, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXFF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXK : CM8INV port map( A => XXDXXXXXXXXXXK, 
                           Y => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXK : CM8INV port map( A => XXDXXXXXXXXXXF, Y
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXDXXXXXYXXXXXXXH : CM8 port map( D0 => axrdata(11), D1 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXX, D3 => axrdata(11),
                           S00 => XXDXXXXDXXXXXYXXXXXXXXXXXXX, S01 => VXXXXXXXX
                           , S10 => axrdata(9), S11 => XXDXXXXXX, Y => 
                           XXDXXXXDXXXXXYXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXL : CM8INV port map( A => XXDXXXXXXXXXXJ, Y
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXYXXXXXXXXXF : XOR4 port map( A => axrdata(3), B => axrdata(11),
                           C => axrdata(7), D => XXDXXXXDXXXXXYXXXXXXXXXXXXXJ, 
                           Y => XXDXXXXDXXXXXYXXXXXH);
   XXDXXXXDXXXXXXFLXXXXXXXX : AND2B port map( A => XXXDXXXXDXXXXYXXXXX, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXX, Y => XXDXXXXXXXXXXFL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => axrdata(16), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D2 => 
                           axrdata(16), D3 => axrdata(16), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXXXXXXXJ, S10 => 
                           XXDXXXXDXXXXXYXXXXXH, S11 => XXDXXXXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXQ);
   XXDXXXXDXXXXXYXXXXXXXJ : CM8 port map( D0 => axrdata(10), D1 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXF, D2 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXF, D3 => axrdata(10)
                           , S00 => XXDXXXXDXXXXXYXXXXXXXXXXXXXF, S01 => 
                           VXXXXXXXX, S10 => axrdata(4), S11 => XXDXXXXXX, Y =>
                           XXDXXXXDXXXXXYXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXL : CM8INV port map( A => XXDXXXXXXXXF, Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXDXXXXXXFLXXXXXXXXF : OR2 port map( A => XXDXXXXDXXXXXYXXXXXK, B => 
                           XXDXXXXDXXXXXYXXXXXL, Y => XXDXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXP : CM8INV port map( A => axrdata(8), Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXQ : CM8INV port map( A => axrdata(9), Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => axrdata(17), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D2 => 
                           axrdata(17), D3 => axrdata(17), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXXXXXXXF, S10 => 
                           XXDXXXXDXXXXXYXXXXXJ, S11 => XXDXXXXDXXXXXXXXF, Y =>
                           XXDXXXXXXXXXXFD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXV : CM8INV port map( A => axrdata(7), Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXW : OR4C port map( A => 
                           XXDXXXXDXXXXXYXXXXXJ, B => XXXDXXXXDXXXXYXXXXX, C =>
                           XXDXXXXDXXXXXYXXXXXH, D => XXDXXXXDXXXXXYXXXXXXXXXXX
                           , Y => XXDXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXP : CM8 port map( D0 => axrdata(2), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D2 => 
                           axrdata(2), D3 => axrdata(2), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXXXXXXXFL, S10 =>
                           XXDXXXXDXXXXXYXXXXXH, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXFQ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXQ : CM8 port map( D0 => axrdata(3), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, D2 => 
                           axrdata(3), D3 => axrdata(3), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXXXXXXXFL, S10 =>
                           XXDXXXXDXXXXXYXXXXXJ, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXHF);
   XXDXXXXDXXXXXYXXXXXXXK : XOR4 port map( A => axrdata(13), B => axrdata(6), C
                           => axrdata(2), D => XXDXXXXDXXXXXYXXXXXXXXXXXXXL, Y 
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXX);
   XXDXXXXDXXXXXYXXXXXXXL : XOR2 port map( A => axrdata(17), B => axrdata(15), 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXFD : CM8INV port map( A => axrdata(6), Y =>
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXP : CM8INV port map( A => axrdata(16), Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXX : OR2B port map( A => XXDXXXXDXXXXXYXXXXXL, 
                           B => XXDXXXXDXXXXXYXXXXXK, Y => XXDXXXXDXXXXXXXXH);
   XXDXXXXDXXXXXYXXXXXXXP : XOR4 port map( A => axrdata(17), B => axrdata(13), 
                           C => axrdata(14), D => axrdata(8), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXX : XOR2 port map( A => XXDXXXXDXXXXXYXXXXXL
                           , B => XXDXXXXDXXXXXXXXXXXXLXXXXXX, Y => 
                           XXXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXX);
   XXDXXXXDXXXXXYXXXXX : CM8 port map( D0 => XXDXXXXDXXXXXYXXXXXXXXXXXXXL, D1 
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXF, D2 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXF, D3 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXL, S00 => 
                           XXDXXXXDXXXXXYXXXXXXXFD, S01 => VXXXXXXXX, S10 => 
                           axrdata(0), S11 => XXDXXXXXX, Y => 
                           XXXDXXXXDXXXXYXXXXX);
   XXDXXXXDXXXXXYXXXXXF : CM8 port map( D0 => XXDXXXXDXXXXXYXXXXXXXXXXXXXK, D1 
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXK, S00 => 
                           XXDXXXXDXXXXXYXXXXXXXFD, S01 => VXXXXXXXX, S10 => 
                           axrdata(1), S11 => XXDXXXXXX, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXK, D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D2 => 
                           XXDXXXXXX, D3 => VXXXXXXXX, S00 => axrdata(15), S01 
                           => VXXXXXXXX, S10 => XXDXXXXDXXXXXXXXH, S11 => 
                           XXDXXXXDXXXXXXXXF, Y => XXDXXXXXXXXXXH);
   XXDXXXXDXXXXXYXXXXXXXQ : XOR2 port map( A => axrdata(16), B => axrdata(14), 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXL : CM8 port map( D0 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, D1 => 
                           XXDXXXXXXXXF, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 
                           => axrdata(14), S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXXXX, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXFV);
   XXDXXXXDXXXXXYXXXXXXXXXXXX : CM8INV port map( A => axrdata(11), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXFF : CM8INV port map( A => axrdata(2), Y =>
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXLXXXXXXXX : XOR4 port map( A => XXDXXXXDXXXXXYXXXXXH, B 
                           => XXDXXXXDXXXXXYXXXXXXXXXXX, C => 
                           XXDXXXXDXXXXXYXXXXXJ, D => XXDXXXXDXXXXXYXXXXXK, Y 
                           => XXDXXXXDXXXXXXXXXXXXLXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : OR2B port map( A => 
                           XXDXXXXDXXXXXYXXXXXH, B => XXDXXXXDXXXXXYXXXXXJ, Y 
                           => XXDXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXQ : CM8INV port map( A => XXDXXXXXXXXF, Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXYXXXXXXXV : XOR2 port map( A => axrdata(9), B => axrdata(7), Y 
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXYXXXXXXXW : XOR2 port map( A => XXDXXXXDXXXXXYXXXXXXXXXXXXXP, B
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXK, Y => 
                           XXDXXXXDXXXXXYXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXFH : CM8INV port map( A => axrdata(3), Y =>
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXV : CM8 port map( D0 => axrdata(6), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, D2 => 
                           axrdata(6), D3 => axrdata(6), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXDXXXXXXXXXX, S10
                           => XXDXXXXDXXXXXYXXXXXH, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXX);
   XXDXXXXDXXXXXYXXXXXXXXXXXXF : CM8INV port map( A => axrdata(10), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXYXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXL, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXW : CM8 port map( D0 => axrdata(7), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, D2 => 
                           axrdata(7), D3 => axrdata(7), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXXXXXXXFL, S10 =>
                           XXDXXXXDXXXXXYXXXXXJ, S11 => XXDXXXXDXXXXXXXXH, Y =>
                           XXDXXXXXXXXXXFJ);
   XXDXXXXDXXXXXYXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXK, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXP : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXDXXXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, S00 => 
                           XXDXXXXXXXXXXJ, S01 => XXDXXXXXXXXXXK, S10 => 
                           axrdata(10), S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXFW)
                           ;
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXX : AND2 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXX, B => XXXDXXXXDXXXXYXXXXX,
                           Y => XXDXXXXDXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXX : OR2A port map( A => XXXDXXXXDXXXXYXXXXX, B 
                           => XXDXXXXDXXXXXYXXXXXXXXXXX, Y => XXDXXXXDXXXXXXXX)
                           ;
   XXDXXXXDXXXXXXFLXXXXXXXXXX : AND2B port map( A => XXDXXXXDXXXXXYXXXXXH, B =>
                           XXDXXXXDXXXXXYXXXXXJ, Y => XXDXXXXXXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXQ : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D2 => 
                           VXXXXXXXX, D3 => XXDXXXXXXXXF, S00 => XXDXXXXXXXXXXF
                           , S01 => XXDXXXXXXXXXXFL, S10 => axrdata(11), S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXF : OR2A port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXX, B => XXXDXXXXDXXXXYXXXXX,
                           Y => XXDXXXXDXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXH, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S10 => 
                           XXDXXXXXXXXXXYXX, S11 => XXDXXXXXXXXXXXXXXXFP, Y => 
                           XXDXXXXXXXXXXYXXF);
   XXDXXXXXXXXXXXXXXXXXXXLXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, D1 => 
                           XXDXXXXXXXXXXXXXXFK, D2 => tmout(19), D3 => 
                           tmout(19), S00 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXW,
                           S01 => XXDXXXXXXXXXXXXXXFW, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => XXDXXXXXX,
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFH);
   XXDXXXXXXXXXXXXXDDXXLX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXJ, D2 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXJ, D3 => XXDXXXXXX, S00
                           => XXDDXXXXXW, S01 => VXXXXXXXX, S10 => XXDDXXXXXV, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXDDXXLXXP);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXX : CM8INV port map( A => axrdata(13), Y => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXF : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXJJ, D1 =>
                           tmout(30), D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP
                           , D3 => tmout(30), S00 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, S11 => 
                           XXDXXXXXXXXXXXXXXXXXV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXK);
   XXDXXXXXXXXXXXXXXX : XOR2 port map( A => XXDDXXXXXF, B => rds(0), Y => 
                           XXDXXXXXXXXXXXXXXXJV);
   XXDXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXXXXXX : AND4 port map( A => XXDDXXXXXK, B => 
                           XXDDXXXXXP, C => XXDDXXXXXJ, D => XXDDXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXWDXXXXXXXX : DFE3C port map( D => XXDXXXXXXXXXXQ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHD, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD);
   XXDXXXXXXXXXXXXXX : OR4 port map( A => XXDXXXXXXXXXXXXXXXXXJ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXHV);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF);
   XXDXXXXXXXXXXXXXXXXXXXXXX : OR4D port map( A => XXDDXXXXXV, B => XXDDXXXXXL,
                           C => XXDDXXXXXW, D => XXDDXXXXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJL);
   XXDXXXXXXXXXXXXXXXXXXXLXXH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, D1 => 
                           XXDXXXXXXXXXXXXXXFW, D2 => tmout(17), D3 => 
                           tmout(17), S00 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFD
                           , S01 => XXDXXXXXXXXXXXXXXFQ, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => XXDXXXXXX,
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXP);
   XXDXXXXXXXXXXXXWDXXXXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXFD, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXDDXXXX : CM8 port map( D0 => VXXXXXXXX, D1 => XXDXXXXXX, D2 
                           => XXDXXXXXX, D3 => VXXXXXXXX, S00 => XXDDXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXXXXXX, S11 => 
                           XXDXXXXXXXXXXYXXXH, Y => XXDXXXXXXXXXXXXXXDDXXXXXFD)
                           ;
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFD, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXP);
   XXDXXXXXXXXXXXXXWDXXXXXXX : CM8 port map( D0 => wdata(0), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXK, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(6));
   XXDXXXXXXXXXXXXXWXDDXXXXX : CM8 port map( D0 => waddr(4), D1 => XXDDXXXXXL, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(4));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXK);
   XXDXXXXXXXXXXXXXXDDXXXXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXV, E
                           => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn, Q
                           => XXDDXXXXXH);
   XXDXXXXXXXXXXXXXDDXXXXXXXXXXX : AND2 port map( A => XXDDXXXXXW, B => 
                           XXDDXXXXXV, Y => XXDXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXDDXXXXXX : CM8 port map( D0 => raddr(11), D1 => XXDDXXXXXX
                           , D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(11));
   XXDXXXXXXXXXXXXXWDXXXXXXXX : CM8 port map( D0 => wdata(8), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXJ, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(14));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXFJ, D1 => 
                           axrdata(7), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rdata(1));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXQ);
   XXDXXXXXXXXXXXXXDDXXLXF : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXX, D2 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10
                           => XXDDXXXXXJ, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXX : AND2A port map( A => 
                           XXDXXXXXXXXXXYXXQ, B => XXXXXXDXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXL, D1 => tmout(39), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D3 => 
                           tmout(39), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, S11 => 
                           XXDXXXXXXXXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXH);
   XXDXXXXXXXXXXXXXDDXX : AND2A port map( A => bypass, B => 
                           XXDXXXXXXXXXXXXXXXHJ, Y => XXDXXXXXXXXXXXXXXDDXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXFF, D3 =>
                           XXDXXXXXX, S00 => XXDXXXXXX, S01 => XXDXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S11 => 
                           XXDXXXXXXXXXXXXXXXHQ, Y => XXDXXXXXXXXXXYXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, D1 => tmout(22)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXP, D3 => 
                           tmout(22), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXFP, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFP);
   XXDXXXXXXXXXXXXX : AND3B port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, 
                           B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, C => 
                           XXDXXXXXXXXXXXXXXFW, Y => XXDXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXDDXXXXX : AND4 port map( A => XXDDXXXXXL, B => XXDDXXXXXK, C
                           => XXDDXXXXXJ, D => XXDDXXXXXH, Y => 
                           XXDXXXXXXXXXXYXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXXF : CM8 port map( D0 => wdata(9), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXP, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(15));
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXHP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXDDXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXF, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXJ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXX, D1 => 
                           axrdata(6), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rdata(0));
   XXDXXXXXXXXXXXXXWXDDXXXXXF : CM8 port map( D0 => waddr(5), D1 => XXDDXXXXXK,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(5));
   XXDXXXXXXXXXXXXXXXDDXXXXXXF : CM8 port map( D0 => raddr(10), D1 => 
                           XXDDXXXXXXF, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10
                           => XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(10));
   XXDXXXXXXXXXXXXXXXXXXXLX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXL, D1 => tmout(6), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, D3 => tmout(6)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXJD, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXP);
   XXDXXXXXXXXXXXXXWDXXXXXXXF : CM8 port map( D0 => wdata(1), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXV, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(7));
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX : AND4A port map( A => XXDXXXXXXXXXXY, B 
                           => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX, C => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXJ, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXX : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXX, S01 => 
                           XXDXXXXXXXXXXYXXV, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXYXXJ);
   XXDXXXXXXXXXXXXXWXDDXXXXXH : CM8 port map( D0 => waddr(8), D1 => XXDDXXXXXF,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(8));
   XXDXXXXXXXXXXXXXXXXXXXLXXL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, D1 => tmout(25)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXV, D3 => 
                           tmout(25), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXJH, S11 
                           => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHK);
   XXDXXXXXXXXXXXXXXXXXXXLXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXW, D1 => tmout(1), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D3 => tmout(1)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ,
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXW);
   XXDXXXXXXXXXXXXXXWXXXXXXXX : AND2B port map( A => re, B => we, Y => 
                           XXDXXXXXXXXXXXXXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXL : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXDDXXXXX : CM8 port map( D0 => raddr(2), D1 => XXDDXXXXXQ, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(2));
   XXDXXXXXXXXXXXXWDXXXXXXX : DFE3C port map( D => XXDXXXXXXXXXXFQ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXWDXXXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXHF, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D1 => XXDXXXXXX, D2
                           => XXDXXXXXXXXXXXXXXXFV, D3 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S00 =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, S01 => 
                           XXXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S11 => 
                           XXXDXXXXDXXXXYXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJF, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXWXDDXXXXXJ : CM8 port map( D0 => waddr(9), D1 => XXDDXXXXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(9));
   XXDXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX : AND4C port map( A => 
                           XXDXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXQXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXX, E => XXDXXXXXXXXXXYXXW,
                           CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXDDXXXXXF : CM8 port map( D0 => raddr(3), D1 => XXDDXXXXXP,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(3));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXH);
   XXDXXXXXXXXXXXXXDDXXLXH : AND2A port map( A => XXDXXXXXXXXXXXXXXXHF, B => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXL);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXV : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXXXXX : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXK, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXL);
   XXDXXXXXXXXXXXXXDDXXXXF : AND2A port map( A => XXYPXXXXXX, B => 
                           XXDXXXXXXXXXXXXXXXHJ, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXW : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFP, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFL, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXXXXXXXXLXH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXQ, D1 => tmout(8), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D3 => tmout(8),
                           S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXHV, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXV);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXH, S00 => 
                           XXDDXXXXXL, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXF, S10 
                           => waddr(4), S11 => XXDXXXXXXXXXXXXXXXHH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXL, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXF : AND3B port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ
                           , B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, C => 
                           XXDXXXXXXXXXXXXXXFQ, Y => XXDXXXXXXXXXXXXXXFW);
   XXDXXXXXXXXXXXXXH : AND3C port map( A => XXDXXXXXXXXXXXXXXXXXV, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, Y => 
                           XXDXXXXXXXXXXXXXXXJJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXXLXXP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXK, D1 => tmout(10), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, D3 => 
                           tmout(10), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01
                           => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXJ, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFV);
   XXDXXXXXXXXXXXXXXXF : OR4 port map( A => XXDXXXXXXXXXXXXXXXXJ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXL : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXV);
   XXDXXXXXXXXXXXXXXXH : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D2 => VXXXXXXXX
                           , D3 => VXXXXXXXX, S00 => XXDXXXXXXXXXXXXXXXXXXXXXXP
                           , S01 => XXDXXXXXXXXXXXXXXFV, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, Y => 
                           XXDXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJJ, D1 => tmout(37), D2 
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXWXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXJP, D1 => 
                           VXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXJP, S00 => XXDDXXXXXX, S01 => 
                           VXXXXXXXX, S10 => waddr(11), S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFW, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFV, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFD : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXQ);
   XXDXXXXXXXXXXXXXWXDDXXXXXK : CM8 port map( D0 => waddr(0), D1 => XXDDXXXXXW,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(0));
   XXDXXXXXXXXXXXXXWXDDXXXXXL : CM8 port map( D0 => waddr(1), D1 => XXDDXXXXXV,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(1));
   XXDXXXXXXXXXXXXXXXXXXXLXXV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, D1 => tmout(18)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXQ, D3 => 
                           tmout(18), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXFW, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFJ);
   XXDXXXXXXXXXXXXXJ : AND3B port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV,
                           B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, C => 
                           XXDXXXXXXXXXXXXXXFP, Y => XXDXXXXXXXXXXXXXXXFW);
   XXDXXXXXXXXXXXXXWDXXXXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXXXXXP, D1 => 
                           wp(3), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXW, D3 => 
                           XXDXXXXXX, S00 => bypass, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S11 => XXDXXXXXX, Y => 
                           axwdata(3));
   XXDXXXXXXXXXXXXXDDXXXXH : AND2A port map( A => XXYPXXXXXX, B => 
                           XXDXXXXXXXXXXXXXXXHJ, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFF);
   XXDXXXXXXXXXXXXXXDDXXXXXH : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXX, E
                           => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn, Q
                           => XXDDXXXXXQ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXFW, D1 => 
                           axrdata(10), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rdata(4));
   XXDXXXXXXXXXXFXXXXLXXD : DFP1B port map( D => XXDXXXXXX, CLK => clk, PRE => 
                           rstn, Q => XXDXXXXXXXXXXXFXXXXLXXDX);
   XXDXXXXXXXXXXXXXWDXXXXXXXXH : CM8 port map( D0 => wdata(5), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXQ, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(11));
   XXDXXXXXXXXXXXXXDDXLDXXXXXXXXXX : AND2 port map( A => XXDXXXXXXXXXXYXXK, B 
                           => XXDXXXXXXXXXXXXXXXDDXX, Y => 
                           XXDXXXXXXXXXXXXXDDXLDXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, D1 => tmout(24)
                           , D2 => XXDXXXXXXXXXXXXXXXJH, D3 => tmout(24), S00 
                           => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXFW, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXQ);
   XXDXXXXXXXXXXXXXWDXXXXXXXXJ : CM8 port map( D0 => wdata(4), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXH, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(10));
   XXDXXXXXXXXXXXXXDDXXLXJ : AND2B port map( A => XXDDXXXXXW, B => 
                           XXDXXXXXXXXXXXXXXXHF, Y => XXDXXXXXXXXXXXXXXDDXXLXXK
                           );
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXYXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXDDXXLXXXXXX : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, Y 
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXFD : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, D1 => tmout(31)
                           , D2 => XXDXXXXXXXXXXXXXXFL, D3 => tmout(31), S00 =>
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXXJJ, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHW);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXJ : CM8 port map( D0 => axrdata(11), D1 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXF, D2 => 
                           axrdata(11), D3 => axrdata(11), S00 => 
                           XXDXXXXXXXXXXF, S01 => XXDXXXXXXXXXXFL, S10 => 
                           bypass, S11 => XXDXXXXXXXXF, Y => rdata(5));
   XXDXXXXXXXXXXXXXXXXXXXLXJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXV, D1 => tmout(0), D2
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => VXXXXXXXX, S10
                           => XXDXXXXXX, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXF);
   XXDXXXXXXXXXXXXXDDXXLXK : CM8 port map( D0 => XXDDXXXXX, D1 => VXXXXXXXX, D2
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => XXDDXXXXXF, 
                           S01 => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXF, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFK, S11 => 
                           XXDXXXXXXXXXXXXXXXHF, Y => XXDXXXXXXXXXXXXXXDDXXLXXJ
                           );
   XXDXXXXXXXXXXXXWDXXXXXXXXH : DFE3C port map( D => XXDXXXXXXXXXXFK, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXWDXXXXXXXJ : CM8 port map( D0 => XXDXXXXXXXXXXXXXXL, D1 => 
                           wp(2), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXJ, D3 => 
                           XXDXXXXXX, S00 => bypass, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S11 => XXDXXXXXX, Y => 
                           axwdata(2));
   XXDXXXXXXXXXXXXXXDDXXXXXJ : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXW, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXP);
   XXDXXXXXXXXXXXXXXXJ : XOR2 port map( A => XXDDXXXXXXF, B => rds(2), Y => 
                           XXDXXXXXXXXXXXXXXXJF);
   XXDXXXXXXXXXXXXPXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXFQ, D1 => 
                           axrdata(2), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rp(2));
   XXDXXXXXXXXXXXXXXXXXXXLXXFF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXF, D1 => tmout(11), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, D3 => 
                           tmout(11), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01
                           => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXK, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFJ, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL);
   XXDXXXXXXXXXXXXXXXK : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, D2 => VXXXXXXXX
                           , D3 => VXXXXXXXX, S00 => XXDXXXXXXXXXXXXXXXXXXXXXXL
                           , S01 => XXDXXXXXXXXXXXXXXXJH, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXF : OR3 port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, B
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXJQ);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXX : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, Y
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFD : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFK, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXFH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D1 => tmout(36),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXJ, D3 => 
                           tmout(36), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXFV, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFQ, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : AND2B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXYXXK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHF, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXP, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXWDXXXXXXXXJ : DFE3C port map( D => XXDXXXXXXXXXXFP, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXXXXW, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXV, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, Y => 
                           XXDXXXXXXXXXXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFH, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXF : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, Y
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXJ);
   XXDXXXXXXXXXXXXLXWDXWXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXXFLXX, E => 
                           XXDXXXXXXXXXXYXXQ, CLK => clk, CLR => rstn, Q => 
                           slowdown);
   XXDXXXXXXXXXXXXPXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXHF, D1 => 
                           axrdata(3), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rp(3));
   XXDXXXXXXXXXXXXXXXXXXXLXK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXK, D1 => tmout(9), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, D3 => tmout(9)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
                           S11 => XXDXXXXXXXXXXXXXXXHV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXX);
   XXDXXXXXXXXXXXXXXWXXXXX : CM8 port map( D0 => waddr(10), D1 => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXXXXX, D2 => VXXXXXXXX, D3 
                           => VXXXXXXXX, S00 => XXDDXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXXHK, S11 => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXX, Y => XXDXXXXXXXXXXY);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXH, D1 
                           => waddr(7), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXDDXXXXXH, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXFQ, S11 => XXDXXXXXXXXXXXXXXXHL, Y
                           => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHH, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXHQ, D2 => XXDXXXXXXXXXXXXXXXXXW, 
                           D3 => XXDXXXXXXXXXXXXXXXXXW, S00 => 
                           XXDXXXXXXXXXXXXXXXDDXX, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXFD, S11 => XXDXXXXXXXXXXXXXXXXXW
                           , Y => XXDXXXXXXXXXXYXXP);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXFLXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXFLXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXL : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, D2 => VXXXXXXXX
                           , D3 => VXXXXXXXX, S00 => XXDXXXXXXXXXXXXXXXXXXXXXXQ
                           , S01 => XXDXXXXXXXXXXXXXXFP, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, Y => 
                           XXDXXXXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXDDXXXXJ : AND4A port map( A => XXDXXXXXXXXXXYXXXH, B => 
                           XXDDXXXXX, C => XXDXXXXXXXXXXYXXX, D => XXDDXXXXXF, 
                           Y => XXDXXXXXXXXXXXXXXDDXXXXXFK);
   XXDXXXXXXXXXXXXXDDXLDXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXYXXK, D1 => 
                           VXXXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXYXXQ, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXXXX, S11 => 
                           XXDXXXXXXXXXXXXXXXHQ, Y => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXX);
   XXDXXXXXXXXXXXXXXXP : XOR2 port map( A => XXDDXXXXX, B => rds(1), Y => 
                           XXDXXXXXXXXXXXXXXXJK);
   XXDXXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXJK, D1 =>
                           VXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXJK, S00 => XXDDXXXXXX, S01 => 
                           VXXXXXXXX, S10 => rds(3), S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJK);
   XXDXXXXXXXXXXXXXXXXXXXLXXFJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, D1 => tmout(16)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, D3 => 
                           tmout(16), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXFQ, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : AND4 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, B => 
                           XXDXXXXXXXXXXXXWXX, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D => 
                           XXDXXXXXXXXXXXXXXDDXXX, Y => XXDXXXXXXXXXXYXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFF, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXJ, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXH : AND2B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, B => 
                           XXDXXXXXXXXXXXXXXXXXFD, Y => XXDXXXXXXXXXXXXXXXJL);
   XXDXXXXXXXXXXXXXXXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXW, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXXDXXXXDXXXXYXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D2 
                           => VXXXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXX, S01 => VXXXXXXXX,
                           S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S11 => 
                           XXDXXXXXXXXXXYXXK, Y => XXDXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXH : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, Y
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXX : DFC1B port map( D => XXDXXXXXXXXXXYXXF, CLK => 
                           clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : OR4 port map( A => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXX, B => 
                           XXDXXXXXXXXXXXXXXXFP, C => XXDXXXXXXXXXXYXX, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXP, D1 => tmout(7), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D3 => tmout(7)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW,
                           S11 => XXDXXXXXXXXXXXXXXXJD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXP);
   XXDXXXXXXXXXXXXXXXQ : XOR2 port map( A => XXDDXXXXXK, B => waddr(5), Y => 
                           XXDXXXXXXXXXXXXXXXHP);
   XXDXXXXXXXXXXXXXDDXXLXL : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXH, D2 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXH, D3 => XXDXXXXXX, S00
                           => XXDDXXXXXJ, S01 => XXDXXXXXXXXXXXXXXDDXXXXXFH, 
                           S10 => XXDDXXXXXH, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXV);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXF);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXXF : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, 
                           Y => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXDXXXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXXJL, E => 
                           XXDXXXXXXXXXXYXXP, CLK => clk, CLR => rstn, Q => 
                           XXXXXXDXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXFK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, D1 => 
                           XXDXXXXXXXXXXXXXXXFW, D2 => tmout(23), D3 => 
                           tmout(23), S00 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXH,
                           S01 => XXDXXXXXXXXXXXXXXFP, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => XXDXXXXXX,
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFW);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXX, D1 => 
                           XXYPXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 =>
                           axrdata(14), S01 => VXXXXXXXX, S10 => XXDXXXXXXXX, 
                           S11 => XXDXXXXXXXXXXXXXXXXXXXXXXXFD, Y => rdata(8));
   XXDXXXXXXXXXXXXXXXDDXXXXXH : CM8 port map( D0 => raddr(7), D1 => XXDDXXXXXH,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(7));
   XXDXXXXXXXXXXXXWDXXXXXXXH : DFE3C port map( D => XXDXXXXXXXXXX, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXWDXXXXXXXJ : DFE3C port map( D => XXDXXXXXXXXXXFJ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXDDXXXXXJ : CM8 port map( D0 => raddr(6), D1 => XXDDXXXXXJ,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(6));
   XXDXXXXXXXXXXXWX : DFC1B port map( D => XXDXXXXXXXXXXYXXL, CLK => clk, CLR 
                           => rstn, Q => XXDXXXXXXXXXXXXWXX);
   XXDXXXXXXXXXXXXXXXXXXXXXF : DFC1B port map( D => XXDXXXXXXXXXXYXXXF, CLK => 
                           clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXL : CM8 port map( D0 => XXDXXXXXXXXXXH, D1 => 
                           axrdata(15), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(9));
   XXDXXXXXXXXXXXXXL : AND4C port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD
                           , B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, D => 
                           XXDXXXXXXXXXXXXXXFP, Y => XXDXXXXXXXXXXXXXXXJH);
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXX : OR3A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXXXXXXXXXXXXXXFD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXFL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, D1 => tmout(38), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, D3 => 
                           tmout(38), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXX, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFW);
   XXDXXXXXXXXXXXXXWDXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXXXXXFD, D1 => 
                           wp(1), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXQ, D3 => 
                           XXDXXXXXX, S00 => bypass, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S11 => XXDXXXXXX, Y => 
                           axwdata(1));
   XXDXXXXXXXXXXXXWDXXXXXXXK : DFE3C port map( D => XXDXXXXXXXXXXFF, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXWXXXXXXXXXX : CM8INV port map( A => waddr(10), Y => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWXDDXXXXXP : CM8 port map( D0 => waddr(3), D1 => XXDDXXXXXP,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(3));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXF);
   XXDXXXXXXXXXXXXXXDDXXXXXK : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXK, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXW);
   XXDXXXXXXXXXXXXXXXDDXXXXXK : CM8 port map( D0 => raddr(9), D1 => XXDDXXXXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(9));
   XXDXXXXXXXXXXXXXWDXXXXXXXXK : CM8 port map( D0 => wdata(7), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXL, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(13));
   XXDXXXXXXXXXXXXXXXXXXXLXXFP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, D1 => tmout(14),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHD, D3 => 
                           tmout(14), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXFH, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXP : CM8 port map( D0 => XXDXXXXXXXXXXFP, D1 => 
                           axrdata(12), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rdata(6));
   XXDXXXXXXXXXXXXXXXXXXXLXXFQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, D1 => tmout(33)
                           , D2 => XXDXXXXXXXXXXXXXXFF, D3 => tmout(33), S00 =>
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXFJ, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXL, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH);
   XXDXXXXXXXXXXXXPXXXXXXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXP, D1 => 
                           axrdata(0), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rp(0));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXX : OR3A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXXXXXXXXXXXXXXFD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX);
   XXDXXXXXXXXXXXXXXDDX : DFE3C port map( D => XXDXXXXXXXXXXXXXXXXXW, E => 
                           XXDXXXXXXXXXXYXXH, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXDDXX);
   XXDXXXXXXXXXXXXXWXDDXXXXXQ : CM8 port map( D0 => waddr(2), D1 => XXDDXXXXXQ,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(2));
   XXDXXXXXXXXXXXXXP : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXXXXQ, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXK, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, Y => 
                           XXDXXXXXXXXXXXXXXFH);
   XXDXXXXXXXXXXXXXWDXXXXXXXXL : CM8 port map( D0 => wdata(6), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXX, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(12));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHF);
   XXDXXXXXXXXXXXXXXXXXXXLXXFV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHH, D1 => tmout(28),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, D3 => 
                           tmout(28), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, S11 => 
                           XXDXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJD);
   XXDXXXXXXXXXXXXXXXDDXXXXXL : CM8 port map( D0 => raddr(8), D1 => XXDDXXXXXF,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(8));
   XXDXXXXXXXXXXXXXXDDXXXXXL : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXP, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXV);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXQ : CM8 port map( D0 => axrdata(13), D1 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXH, D2 => 
                           axrdata(13), D3 => axrdata(13), S00 => 
                           XXDXXXXXXXXXXJ, S01 => XXDXXXXXXXXXXFL, S10 => 
                           XXYPXXXXXX, S11 => XXDXXXXXXXXF, Y => rdata(7));
   XXDXXXXXXXXXXXXXWDXXXXXXXL : CM8 port map( D0 => XXDXXXXXXXXXXXXXXW, D1 => 
                           wp(0), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXX, D3 => 
                           XXDXXXXXX, S00 => bypass, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S11 => XXDXXXXXX, Y => 
                           axwdata(0));
   XXDXXXXXXXXXXXXWDXXXXXXXL : DFE3C port map( D => XXDXXXXXXXXXXW, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXV : XOR2 port map( A => XXDDXXXXXQ, B => waddr(2), Y => 
                           XXDXXXXXXXXXXXXXXXHL);
   XXDXXXXXXXXXXXXWDXXXXXXXXK : DFE3C port map( D => XXDXXXXXXXXXXV, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXX, D1 => 
                           VXXXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXYXXQ, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, S11 => 
                           XXDXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXX, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXHH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXK, E => XXDXXXXXXXXXXYXXW
                           , CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXXXXXXYXXV, D3 => XXDXXXXXX,
                           S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S01 
                           => VXXXXXXXX, S10 => XXDXXXXXXXXXXYXXK, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXYXXXF);
   XXDXXXXXXXXXXXXXXXFLXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXFLXXXXXXXXXXXXX, D1 => XXDXXXXXX,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXH, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, S11 => 
                           XXXXXXDXXXX, Y => XXDXXXXXXXXXXXXXXXFLXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHW, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF);
   XXDXXXXXXXXXXXXXXH : OR3 port map( A => XXDXXXXXXXXXXXXXXXHV, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => XXDXXXXXXXXXXXXXXXJF, 
                           Y => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXWDXXXXXXXP : DFE3C port map( D => XXDXXXXXXXXXXL, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXLXXFW : CM8 port map( D0 => XXDXXXXXXXXXXXXXXFH, D1 =>
                           tmout(13), D2 => XXDXXXXXXXXXXXXXXXXF, D3 => 
                           tmout(13), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJK, D2 => VXXXXXXXX, D3 
                           => VXXXXXXXX, S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXJ
                           , S01 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXJV, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJL, Y => 
                           XXDXXXXXXXXXXXXXXXHQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXV, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHD : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJD, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH);
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXHQ, D2 => XXDXXXXXXXXXXXXXXXXXW, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXXDDXX, S01 
                           => XXDXXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S11 => 
                           XXDXXXXXXXXXXXXXXXXXFD, Y => XXDXXXXXXXXXXYXXH);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D2 => VXXXXXXXX, D3
                           => VXXXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXX, S01 => 
                           XXDXXXXXXXXXXXXXXXHD, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, S11 => XXDXXXXXX, Y
                           => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXLXP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXX, D1 => tmout(5), D2 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D3 => tmout(5)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXJ, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXQ);
   XXDXXXXXXXXXXXXXDDXXLXP : CM8 port map( D0 => XXDDXXXXXK, D1 => VXXXXXXXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => XXDDXXXXXL,
                           S01 => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXK, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S11 => 
                           XXDXXXXXXXXXXXXXXXHF, Y => XXDXXXXXXXXXXXXXXDDXXLXXQ
                           );
   XXDXXXXXXXXXXXXXXXXXXXLXXHD : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, D1 => 
                           XXDXXXXXXXXXXXXXXFP, D2 => tmout(21), D3 => 
                           tmout(21), S00 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFP
                           , S01 => XXDXXXXXXXXXXXXXXFK, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => XXDXXXXXX,
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHV);
   XXDXXXXXXXXXXXXWDXXXXXXXXL : DFE3C port map( D => XXDXXXXXXXXXXFW, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXXXXXP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXQ, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFL : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHH);
   XXDXXXXXXXXXXXXPXXXXXXXXXJ : CM8 port map( D0 => XXDXXXXXXXXXXFH, D1 => 
                           axrdata(1), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rp(1));
   XXDXXXXXXXXXXXXXXXW : XOR2 port map( A => XXDDXXXXXF, B => waddr(8), Y => 
                           XXDXXXXXXXXXXXXXXXHK);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXX, D1 => 
                           VXXXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXFD, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, S11 => 
                           XXDXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXQ : DFE3C port map( D => XXDXXXXXXXXXXXXXXXHW, E => 
                           XXDXXXXXXXXXXYXXJ, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXHD);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXX : AND2A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXFD, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXDDXXLXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXXF, D2 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXXF, D3 => XXDXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXDDXXXXXFK, S01 => VXXXXXXXX,
                           S10 => XXDDXXXXXXF, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXDXXXXX : AND2 port map( A => XXDXXXXXXXXXXXXWXX, 
                           B => XXDXXXXXXXXXXXXXXDDXXXXXFF, Y => 
                           scrub_corrected);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXV : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXH, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHJ, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHK, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXLXQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXJ, D1 => tmout(2), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D3 => 
                           tmout(2), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 
                           => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXK);
   XXDXXXXXXXXXXXXXDDXLDXXX : CM8 port map( D0 => VXXXXXXXX, D1 => XXDXXXXXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXDDXLDXXXXXXXX, S01 => 
                           XXDXXXXXXXXXXYXXV, S10 => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXX, S11 => XXDXXXXXX, Y =>
                           XXDXXXXXXXXXXXXXDDXXF);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXX : OR2 port map( A => 
                           XXDXXXXXXXXXXXFXXXXLXXDX, B => stop_scrub, Y => 
                           XXDXXXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXLXXHF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFV, D1 => tmout(26),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, D3 => 
                           tmout(26), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXQ, S11 
                           => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFF);
   XXDXXXXXXXXXXXXXV : AND3B port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV
                           , B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, C => 
                           XXDXXXXXXXXXXXXXXFK, Y => XXDXXXXXXXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXL);
   XXDXXXXXXXXXXXXXDDXXLXQ : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXQ, D2 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXQ, D3 => XXDXXXXXX, S00
                           => XXDXXXXXXXXXXXXXXXXXL, S01 => VXXXXXXXX, S10 => 
                           XXDDXXXXXQ, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXX);
   XXDXXXXXXXXXXXXXDDXXXXXF : NAND4 port map( A => XXDDXXXXXW, B => XXDDXXXXXV,
                           C => XXDDXXXXXQ, D => XXDDXXXXXP, Y => 
                           XXDXXXXXXXXXXYXXXH);
   XXDXXXXXXXXXXXXXXXFD : OR4A port map( A => XXDXXXXXXXXXXXXXXXFW, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFV : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXQ, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXXDXXXXDXXXXYXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXWXXXXXX : CM8 port map( D0 => we, D1 => XXDXXXXXXXXXXXXWXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFF, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwe);
   XXDXXXXXXXXXXXXXW : AND4C port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK
                           , B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, D => 
                           XXDXXXXXXXXXXXXXXXJJ, Y => XXDXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXW : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXH);
   XXDXXXXXXXXXXXXXDDXXXXK : AND2A port map( A => XXYPXXXXXX, B => 
                           XXDXXXXXXXXXXXXXXXHJ, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXP, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF, S00 => 
                           XXDDXXXXXJ, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXX, S10 
                           => waddr(6), S11 => XXDXXXXXXXXXXXXXXXHP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXHH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHJ, D1 => tmout(41),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, D3 => 
                           tmout(41), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, S11 => 
                           XXDXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXX);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => 
                           waddr(7), Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFW : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXX : OR2A port map( A => XXDXXXXXXXXXXXXXXXHQ, B => 
                           XXDXXXXXXXXXXYXXQ, Y => XXDXXXXXXXXXXXXXXXHF);
   XXDXXXXXXXXXXXXWDXXXXXXXQ : DFE3C port map( D => XXDXXXXXXXXXXHD, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXQ, D1 => 
                           axrdata(16), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(10));
   XXDXXXXXXXXXXXXXXXDDXXXXXP : CM8 port map( D0 => raddr(5), D1 => XXDDXXXXXK,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(5));
   XXDXXXXXXXXXXXXXXXXXXXLXXHJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, D1 => tmout(34)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFK, D3 => 
                           tmout(34), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXFF, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXV);
   XXDXXXXXXXXXXXXXXXXXXLDXXXXXXXX : AND2A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXFD, B => XXDXXXXXXXXXXXXXXXFLXX,
                           Y => XXDXXXXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXXXXDDXXXXXQ : CM8 port map( D0 => raddr(4), D1 => XXDDXXXXXL,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(4));
   XXDXXXXXXXXXXXXXDDXXLXV : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXP, D2 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXP, D3 => XXDXXXXXX, S00
                           => XXDDXXXXXQ, S01 => XXDXXXXXXXXXXXXXXXXXL, S10 => 
                           XXDDXXXXXP, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXW);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXFD, D1 => 
                           axrdata(17), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(11));
   XXDXXXXXXXXXXXXXXJ : OR3 port map( A => XXDXXXXXXXXXXXXXXXJQ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXL : AND2A port map( A => XXDXXXXXXXXXXYXXQ, B => 
                           XXDXXXXXXXXXXYXXK, Y => XXDXXXXXXXXXXXXXXXHW);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHD : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFH);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFQ);
   XXDXXXXXXXXXXXXXXXFF : XOR2 port map( A => XXDDXXXXXW, B => waddr(0), Y => 
                           XXDXXXXXXXXXXXXXXXHH);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXJ);
   XXDXXXXXXXXXXXXXDDXXXXL : AND3A port map( A => XXDXXXXXXXXXXYXXXH, B => 
                           XXDDXXXXXK, C => XXDDXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH);
   XXDXXXXXXXXXXXXWDXXXXXXXXP : DFE3C port map( D => XXDXXXXXXXXXXFV, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXK : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, Y
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXL);
   XXDXXXXXXXXXXXXPXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXL, D1 => 
                           axrdata(5), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rp(5));
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX : OR2 port map( A => 
                           XXDXXXXXXXXXXXFXXXXLXXDX, B => stop_scrub, Y => 
                           XXDXXXXXXXXXXYXXQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : AND4A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXXXXXXXXXXXXHD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXFV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHL, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP);
   XXDXXXXXXXXXXXXXXDDXXXXXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXXF,
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXX);
   XXDXXXXXXXXXXXXXXK : OR4 port map( A => XXDXXXXXXXXXXXXXXXJQ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXXXXXXXXXXXXJD);
   XXDXXXXXXXXXXXXXXDDXXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXX,
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXV, E => XXDXXXXXXXXXXYXXW
                           , CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXHK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFW, D1 => tmout(27),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D3 => 
                           tmout(27), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXK, S11 
                           => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHH);
   XXDXXXXXXXXXXXXXXXXXXLDXXXXXX : AND2A port map( A => XXDXXXXXXXXXXYXXQ, B =>
                           XXDXXXXXXXXXXXXXXXFLXX, Y => XXDXXXXXXXXXXYXXW);
   XXDXXXXXXXXXXXXXXXXXXXLXV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXH, D1 => tmout(3), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, D3 => tmout(3)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXJQ, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXL);
   XXDXXXXXXXXXXXXWDXXXXXXXXQ : DFE3C port map( D => XXDXXXXXXXXXXH, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXFH : XOR2 port map( A => XXDDXXXXX, B => waddr(9), Y => 
                           XXDXXXXXXXXXXXXXXXJP);
   XXDXXXXXXXXXXXXPXXXXXXXXXL : CM8 port map( D0 => XXDXXXXXXXXXXHD, D1 => 
                           axrdata(4), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rp(4));
   XXDXXXXXXXXXXXXXXXFJ : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, D2 => VXXXXXXXX
                           , D3 => VXXXXXXXX, S00 => XXDXXXXXXXXXXXXXXXXXXXXXXK
                           , S01 => XXDXXXXXXXXXXXXXXFF, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXX : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXY, D2 => XXDXXXXXX, D3 => XXDXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX, S01
                           => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXJ, S10 =>
                           XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXYXXL);
   XXDXXXXXXXXXXXXXWXDDXXXXXV : CM8 port map( D0 => waddr(6), D1 => XXDDXXXXXJ,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(6));
   XXDXXXXXXXXXXXXXXXXXXXLXXHL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH, D1 => 
                           XXDXXXXXXXXXXXXXXFQ, D2 => tmout(15), D3 => 
                           tmout(15), S00 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHF
                           , S01 => XXDXXXXXXXXXXXXXXFH, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => XXDXXXXXX,
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXP : CM8 port map( D0 => XXDXXXXXXXXXXXXXXV, D1 => 
                           wp(4), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXF, D3 => 
                           XXDXXXXXX, S00 => bypass, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S11 => XXDXXXXXX, Y => 
                           axwdata(4));
   XXDXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJP);
   XXDXXXXXXXXXXXXXXDDXXXXXP : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXQ, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXFK : XOR2 port map( A => XXDDXXXXXV, B => waddr(1), Y => 
                           XXDXXXXXXXXXXXXXXXFQ);
   XXDXXXXXXXXXXXXXXDDXXXXXQ : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXJ, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXX);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXV : CM8 port map( D0 => XXDXXXXXXXXXXFF, D1 => 
                           axrdata(8), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rdata(2));
   XXDXXXXXXXXXXXXXXXXXXXLXXHP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFH, D1 => tmout(12),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, D3 => 
                           tmout(12), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S11 => 
                           XXDXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHQ);
   XXDXXXXXXXXXXXXXXXXXXLDXXXXXXXXF : AND2A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXFD, B => XXDXXXXXXXXXXXXXXXFLXX,
                           Y => XXDXXXXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXWXDDXXXXXX : CM8 port map( D0 => waddr(10), D1 => 
                           XXDDXXXXXXF, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFL, S01 => VXXXXXXXX, S10
                           => XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(10));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXW : CM8 port map( D0 => XXDXXXXXXXXXXW, D1 => 
                           axrdata(9), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rdata(3));
   XXDXXXXXXXXXXXXXWDXXXXXXXXP : CM8 port map( D0 => wdata(10), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXF, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(16));
   XXDXXXXXXXXXXXXXXXXXXXLXXHQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP, D1 => 
                           XXDXXXXXXXXXXXXXXFV, D2 => tmout(35), D3 => 
                           tmout(35), S00 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFL
                           , S01 => XXDXXXXXXXXXXXXXXFF, S10 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S11 => XXDXXXXXX, 
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHL);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXL : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, Y
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXQ);
   XXDXXXXXXXXXXXXXFD : AND3B port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ
                           , B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, C => 
                           XXDXXXXXXXXXXXXXXXJJ, Y => XXDXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXFF : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXXXXV, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXF, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH, Y => 
                           XXDXXXXXXXXXXXXXXFQ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXF : CM8INV port map( A => axrdata(11), Y =>
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXXQ : CM8 port map( D0 => wdata(11), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXK, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(17));
   XXDXXXXXXXXXXXXXXXXXXXLXXHV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHK, D1 => tmout(40),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, D3 => 
                           tmout(40), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXH, S11 
                           => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXJF);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHK);
   XXDXXXXXXXXXXXXXWXDDXXXXXW : CM8 port map( D0 => waddr(7), D1 => XXDDXXXXXH,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(7));
   XXDXXXXXXXXXXXXXWDXXXXXXXQ : CM8 port map( D0 => XXDXXXXXXXXXXXXXXQ, D1 => 
                           wp(5), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXP, D3 => 
                           XXDXXXXXX, S00 => bypass, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S11 => XXDXXXXXX, Y => 
                           axwdata(5));
   XXDXXXXXXXXXXXXXWXDDXXXXXXF : CM8 port map( D0 => waddr(11), D1 => 
                           XXDDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXDXXXXXXXXXXXXXXDDXXXXXFL, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(11));
   XXDXXXXXXXXXXXXXFH : AND4C port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, D => 
                           XXDXXXXXXXXXXXXXXFJ, Y => XXDXXXXXXXXXXXXXXFV);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => we, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           we, S01 => XXDDXXXXXP, S10 => waddr(3), S11 => 
                           XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXH : CM8INV port map( A => XXYPXXXXXX, Y => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXDDXXXXXV : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXH, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXL);
   XXDXXXXXXXXXXXXXXXXFLXX : DFC1B port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => tmoutflg);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXP : CM8INV port map( A => XXDXXXXXXXXXXYXXXH, Y 
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXX : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXXXXXXXXXXXHQ, D3 => 
                           XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXDDXX, S11
                           => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXDDXLDXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXDDXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXXLXXHW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFQ, D1 => tmout(29),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, D3 => 
                           tmout(29), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXV, S11 
                           => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXL);
   XXDXXXXXXXXXXXXXWDXXXXXXXV : CM8 port map( D0 => wdata(2), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXL, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(8));
   XXDXXXXXXXXXXXXXXXDDXXXXXV : CM8 port map( D0 => raddr(0), D1 => XXDDXXXXXW,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(0));
   XXDXXXXXXXXXXXXWDXXXXXXXV : DFE3C port map( D => XXDXXXXXXXXXXFH, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D1 => VXXXXXXXX, D2
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => XXDXXXXXXXXXXXXXXXHD,
                           S10 => XXDXXXXXXXXXXYXXK, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXDDXXXXXXXXX : CM8INV port map( A => XXDXXXXXXXXXXYXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXW : CM8 port map( D0 => wdata(3), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXH, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(9));
   XXDXXXXXXXXXXXXWDXXXXXXXW : DFE3C port map( D => XXDXXXXXXXXXXP, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXJD : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, D1 => tmout(32),
                           D2 => XXDXXXXXXXXXXXXXXFJ, D3 => tmout(32), S00 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXFL, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFK);
   XXDXXXXXXXXXXXXXXDDXXXXXW : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXL, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXF);
   XXDXXXXXXXXXXXXXXXDDXXXXXW : CM8 port map( D0 => raddr(1), D1 => XXDDXXXXXV,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(1));
   XXDXXXXXXXXXXXXXXXXXXXLXW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXF, D1 => tmout(4), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, D3 => tmout(4)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK,
                           S11 => XXDXXXXXXXXXXXXXXXJQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXH);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXH, E => XXDXXXXXXXXXXYXXW
                           , CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJ, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV);
   XXDXXXXXXXXXXXXXDDXXLXXF : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXX, D2 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXX, D3 => XXDXXXXXX, S00
                           => XXDDXXXXXXF, S01 => XXDXXXXXXXXXXXXXXDDXXXXXFK, 
                           S10 => XXDDXXXXXX, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXF, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXF, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW);
   XXDXXXXXXXXXXXXXXXFL : OR4 port map( A => XXDXXXXXXXXXXXXXXXHV, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, Y => 
                           XXDXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXXXXXXXF, D1 => 
                           VXXXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXFD, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, S11 => 
                           XXDXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXF : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => VXXXXXXXX, D3 => XXDXXXXXXXXXXXXWXX
                           , S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXDDXXX, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXQ : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHF, Y
                           => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXF : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXX, D2 => 
                           VXXXXXXXX, D3 => XXDXXXXXX, S00 => XXXXXXDXXXX, S01 
                           => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, S11 => 
                           XXDXXXXXXXXXXXXXXXXH, Y => XXDXXXXXXXXXXYXXV);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXF : OR3 port map( A => XXDXXXXXXXXXXXXXXXFP
                           , B => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXF, C => 
                           XXDXXXXXXXXXXYXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJD : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHP, E => 
                           XXDXXXXXXXXXXYXXW, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK);
   XXDXXXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => XXDXXXXXX, D1 => VXXXXXXXX,
                           D2 => VXXXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, S01 => 
                           XXDXXXXXXXXXXXXXXFV, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXXXXXJJ);
   XXDXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => re, D1 => XXDXXXXXXXXXXXXXXXHD,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFF, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axre);
   XXDXXXXXXXXXXXXXDDXXLXW : CM8 port map( D0 => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXL
                           , D1 => XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXL, S00 => 
                           XXDXXXXXXXXXXYXXXH, S01 => VXXXXXXXX, S10 => 
                           XXDDXXXXXL, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXJF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, D1 => tmout(20)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFJ, D3 => 
                           tmout(20), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXFK, S11 =>
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXW, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHQ, E => 
                           XXDXXXXXXXXXXXXXXXXXP, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXDDXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHV, E => 
                           XXDXXXXXXXXXXXXXXXXXFF, CLK => clk, CLR => rstn, Q 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV);
   XXDXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => VXXXXXXXX, D1 => VXXXXXXXX, D2 
                           => XXDXXXXXX, D3 => XXDXXXXXXXXXXFL, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJP, S01 => XXDXXXXXXXXXXK
                           , S10 => stop_scrub, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXXDXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXH : DFC1B port map( D => XXDXXXXXXXXXXYXXXJ, CLK => 
                           clk, CLR => rstn, Q => XXDXXXXXXXXXXXXXXXXXXXXXXXFF)
                           ;
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHJ);

end SYN_DEF_ARCH;
