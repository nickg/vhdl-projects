use WORK.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use Std.TextIO.all;
use work.debugtools.all;

ENTITY ram8x32k IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    clkb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ram8x32k;

architecture behavioural of ram8x32k is

  type ram_t is array (0 to 32767) of std_logic_vector(7 downto 0);
  shared variable ram : ram_t := (x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"36",x"35",x"55",x"43",x"4F",x"4E",x"46",x"49",x"47",x"55",x"52",x"45",x"20",x"4D",x"45",x"47",x"41",x"36",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B4",x"1A",x"0D",x"08",x"50",x"08",x"30",x"23",x"01",x"08",x"0B",x"08",x"37",x"01",x"9E",x"32",x"30",x"36",x"31",x"00",x"00",x"00",x"BA",x"BD",x"B6",x"21",x"9D",x"FC",x"00",x"CA",x"D0",x"F7",x"A0",x"35",x"4C",x"68",x"21",x"20",x"81",x"06",x"58",x"9C",x"D5",x"E0",x"37",x"0B",x"5A",x"0C",x"56",x"2A",x"05",x"AB",x"92",x"03",x"D2",x"F4",x"89",x"7E",x"0E",x"A4",x"01",x"0F",x"04",x"00",x"DF",x"63",x"C0",x"DE",x"02",x"20",x"2C",x"D8",x"DB",x"DD",x"E6",x"76",x"DB",x"03",x"0F",x"02",x"02",x"3D",x"AD",x"F3",x"2F",x"F6",x"76",x"B7",x"B9",x"DD",x"F6",x"0C",x"80",x"0A",x"B5",x"07",x"0D",x"56",x"0E",x"A0",x"30",x"E2",x"EF",x"4E",x"CA",x"A8",x"70",x"F2",x"A6",x"99",x"3B",x"EE",x"31",x"8B",x"DD",x"63",x"D5",x"EA",x"6F",x"A6",x"6B",x"DA",x"B4",x"E0",x"B0",x"00",x"4C",x"00",x"5D",x"42",x"2F",x"0D",x"CD",x"4D",x"73",x"41",x"BE",x"9C",x"0A",x"31",x"2E",x"D1",x"30",x"15",x"90",x"40",x"4F",x"F4",x"39",x"18",x"A3",x"46",x"A4",x"24",x"6A",x"30",x"67",x"2D",x"8E",x"39",x"18",x"B4",x"40",x"D1",x"2F",x"08",x"95",x"DA",x"1A",x"80",x"5C",x"42",x"27",x"45",x"D7",x"63",x"09",x"D0",x"00",x"E5",x"19",x"C0",x"45",x"0F",x"E2",x"A2",x"3F",x"1C",x"C0",x"B0",x"B7",x"02",x"D0",x"37",x"05",x"17",x"56",x"CC",x"E5",x"3E",x"D8",x"79",x"97",x"6C",x"36",x"EA",x"50",x"3F",x"1D",x"61",x"27",x"06",x"D6",x"64",x"74",x"E3",x"44",x"7C",x"33",x"B1",x"12",x"0C",x"77",x"22",x"8D",x"45",x"71",x"B9",x"1B",x"E8",x"19",x"BF",x"4C",x"3F",x"19",x"F0",x"24",x"13",x"61",x"84",x"6E",x"07",x"3F",x"16",x"BE",x"1A",x"70",x"3C",x"90",x"98",x"97",x"D7",x"74",x"D2",x"CE",x"7B",x"12",x"80",x"3A",x"86",x"02",x"42",x"95",x"BC",x"D8",x"06",x"77",x"24",x"DA",x"29",x"9D",x"8A",x"20",x"83",x"8E",x"64",x"D5",x"1F",x"5A",x"B6",x"80",x"9A",x"6C",x"0D",x"8D",x"1B",x"21",x"26",x"03",x"28",x"6E",x"97",x"4E",x"71",x"4B",x"22",x"1C",x"55",x"D9",x"3A",x"D9",x"46",x"A0",x"71",x"B1",x"C5",x"14",x"61",x"19",x"66",x"31",x"CD",x"33",x"B4",x"0E",x"26",x"9E",x"90",x"AC",x"66",x"1D",x"2F",x"25",x"B5",x"67",x"45",x"A5",x"2E",x"25",x"65",x"DE",x"ED",x"A6",x"D1",x"22",x"A3",x"64",x"92",x"12",x"B2",x"32",x"92",x"6A",x"68",x"C5",x"39",x"CE",x"09",x"A3",x"1C",x"93",x"32",x"2F",x"66",x"E8",x"34",x"A7",x"E2",x"60",x"8E",x"29",x"62",x"9B",x"77",x"5A",x"D0",x"D4",x"0A",x"D1",x"26",x"B0",x"8A",x"63",x"C1",x"D0",x"72",x"53",x"BE",x"70",x"2F",x"1D",x"B2",x"77",x"C5",x"22",x"2C",x"1C",x"16",x"17",x"BF",x"B2",x"20",x"21",x"29",x"69",x"6C",x"0B",x"9A",x"70",x"05",x"82",x"0C",x"B3",x"A3",x"64",x"73",x"FC",x"63",x"B4",x"32",x"12",x"0C",x"97",x"6E",x"A7",x"C3",x"40",x"2E",x"23",x"F1",x"38",x"63",x"4D",x"79",x"A4",x"68",x"9D",x"91",x"B5",x"62",x"BC",x"E5",x"B4",x"43",x"9D",x"6C",x"D1",x"B2",x"17",x"92",x"D0",x"62",x"2A",x"2C",x"B5",x"29",x"80",x"17",x"EE",x"17",x"47",x"2E",x"24",x"34",x"4B",x"72",x"D5",x"FA",x"56",x"A2",x"10",x"1C",x"32",x"07",x"C6",x"85",x"D0",x"5D",x"E5",x"B5",x"38",x"79",x"2E",x"A7",x"C2",x"2A",x"21",x"63",x"14",x"29",x"10",x"23",x"90",x"85",x"4A",x"1F",x"13",x"6B",x"5B",x"06",x"BE",x"72",x"0A",x"17",x"75",x"32",x"0C",x"BD",x"77",x"D6",x"EB",x"46",x"64",x"B5",x"73",x"2C",x"A3",x"9E",x"52",x"3D",x"10",x"48",x"99",x"BA",x"40",x"DC",x"37",x"00",x"85",x"7D",x"82",x"66",x"CC",x"6A",x"E6",x"0A",x"68",x"51",x"22",x"2D",x"83",x"54",x"76",x"D6",x"83",x"59",x"A7",x"0B",x"BF",x"32",x"E4",x"0B",x"B4",x"CA",x"06",x"16",x"D0",x"22",x"B6",x"C6",x"C1",x"91",x"66",x"72",x"67",x"75",x"5A",x"41",x"A1",x"2B",x"A0",x"56",x"6F",x"4A",x"DC",x"B4",x"38",x"21",x"24",x"D1",x"36",x"59",x"C9",x"77",x"3E",x"6C",x"9D",x"A5",x"51",x"4E",x"6D",x"49",x"39",x"AC",x"1B",x"68",x"CD",x"A7",x"10",x"83",x"A3",x"72",x"43",x"CF",x"D0",x"B8",x"9B",x"27",x"1A",x"21",x"D5",x"09",x"4E",x"8F",x"6D",x"BC",x"74",x"B3",x"B1",x"B1",x"15",x"A0",x"73",x"17",x"16",x"71",x"75",x"69",x"FB",x"A4",x"49",x"66",x"29",x"92",x"68",x"5B",x"02",x"D1",x"2E",x"1F",x"C3",x"70",x"19",x"61",x"B6",x"73",x"03",x"DC",x"D9",x"DC",x"BA",x"38",x"79",x"15",x"5B",x"72",x"3B",x"ED",x"5C",x"E7",x"AF",x"CE",x"CF",x"88",x"1E",x"53",x"DB",x"24",x"91",x"19",x"3A",x"EA",x"8D",x"58",x"64",x"C7",x"24",x"DA",x"EB",x"21",x"F8",x"75",x"65",x"2E",x"FB",x"4C",x"B0",x"07",x"6F",x"63",x"94",x"0D",x"64",x"A5",x"D8",x"C5",x"5A",x"26",x"DD",x"6B",x"FD",x"0C",x"00",x"E8",x"09",x"FF",x"08",x"20",x"40",x"34",x"01",x"1B",x"31",x"4C",x"00",x"04",x"36",x"31",x"58",x"E0",x"01",x"B8",x"02",x"16",x"CA",x"57",x"07",x"5D",x"42",x"4E",x"06",x"6E",x"C7",x"C8",x"9E",x"44",x"6D",x"15",x"4B",x"24",x"A1",x"70",x"44",x"33",x"35",x"1F",x"3C",x"85",x"0A",x"17",x"05",x"00",x"08",x"EF",x"21",x"6A",x"6F",x"79",x"6F",x"EF",x"33",x"76",x"F7",x"32",x"5A",x"FB",x"C6",x"DF",x"61",x"36",x"A0",x"75",x"D2",x"5C",x"1A",x"A7",x"72",x"28",x"B7",x"1A",x"0C",x"31",x"73",x"94",x"E2",x"6E",x"44",x"38",x"43",x"0A",x"6A",x"67",x"0C",x"5A",x"16",x"30",x"00",x"61",x"FA",x"E6",x"6F",x"F0",x"0F",x"74",x"ED",x"B5",x"B3",x"09",x"68",x"50",x"11",x"6D",x"BA",x"23",x"5F",x"CE",x"70",x"F3",x"01",x"78",x"B7",x"BB",x"B7",x"65",x"0D",x"A5",x"9C",x"6F",x"04",x"6D",x"2D",x"6C",x"80",x"79",x"8C",x"78",x"24",x"8A",x"55",x"62",x"64",x"25",x"B8",x"8C",x"63",x"0D",x"B2",x"76",x"04",x"5C",x"43",x"13",x"89",x"33",x"82",x"DC",x"ED",x"6D",x"D9",x"3C",x"A0",x"72",x"7F",x"2A",x"35",x"32",x"D4",x"33",x"29",x"05",x"2F",x"38",x"62",x"72",x"04",x"0D",x"F7",x"15",x"66",x"A9",x"76",x"9F",x"1B",x"E1",x"35",x"42",x"76",x"6F",x"A2",x"40",x"6C",x"AB",x"2A",x"11",x"55",x"63",x"A3",x"DA",x"0D",x"D2",x"11",x"33",x"C1",x"2E",x"35",x"22",x"9F",x"5C",x"E3",x"2A",x"E7",x"D9",x"6C",x"8C",x"CE",x"30",x"6D",x"00",x"35",x"50",x"1F",x"65",x"07",x"E9",x"2B",x"6B",x"20",x"1B",x"61",x"67",x"EE",x"A5",x"03",x"2C",x"20",x"0F",x"AA",x"8B",x"1F",x"6C",x"9B",x"1C",x"E5",x"13",x"66",x"6E",x"6D",x"69",x"75",x"0B",x"4A",x"6F",x"EA",x"A2",x"28",x"E4",x"B7",x"70",x"CD",x"78",x"4C",x"6D",x"AB",x"9D",x"29",x"3A",x"CB",x"07",x"87",x"73",x"5A",x"03",x"06",x"51",x"E9",x"61",x"62",x"6C",x"DE",x"92",x"50",x"0E",x"02",x"AE",x"A1",x"0B",x"B6",x"5F",x"63",x"65",x"EF",x"1E",x"3A",x"13",x"70",x"F7",x"A7",x"48",x"AB",x"99",x"35",x"82",x"37",x"53",x"92",x"6E",x"36",x"DC",x"03",x"B4",x"36",x"45",x"68",x"7A",x"BD",x"37",x"B7",x"32",x"47",x"2A",x"34",x"B3",x"3B",x"C9",x"0D",x"00",x"02",x"0E",x"7D",x"9D",x"67",x"A5",x"0D",x"65",x"20",x"3B",x"B7",x"96",x"D5",x"3A",x"15",x"3D",x"89",x"58",x"35",x"15",x"AB",x"D9",x"8A",x"29",x"66",x"13",x"86",x"64",x"11",x"3D",x"79",x"6C",x"4A",x"4B",x"28",x"DB",x"B0",x"1C",x"19",x"29",x"21",x"AB",x"D3",x"0E",x"63",x"72",x"7D",x"E4",x"65",x"6D",x"5D",x"E8",x"6D",x"8D",x"05",x"0B",x"4C",x"0F",x"DE",x"40",x"0D",x"CA",x"EC",x"04",x"41",x"70",x"CA",x"82",x"3A",x"06",x"B7",x"94",x"04",x"6D",x"70",x"6C",x"83",x"22",x"96",x"72",x"0F",x"73",x"AF",x"36",x"67",x"B6",x"21",x"D4",x"DC",x"61",x"74",x"66",x"6E",x"3A",x"DC",x"36",x"55",x"31",x"04",x"EC",x"35",x"38",x"D0",x"30",x"81",x"32",x"15",x"2A",x"77",x"DA",x"70",x"14",x"B5",x"ED",x"F8",x"96",x"82",x"63",x"68",x"DB",x"EF",x"6E",x"6C",x"AA",x"49",x"02",x"6E",x"F7",x"4B",x"79",x"14",x"E8",x"78",x"01",x"10",x"32",x"B4",x"73",x"77",x"2E",x"B8",x"6D",x"70",x"6C",x"3D",x"84",x"69",x"65",x"72",x"3A",x"DC",x"46",x"66",x"A0",x"02",x"AB",x"9D",x"A8",x"D4",x"00",x"80",x"0E",x"64",x"7B",x"1F",x"6C",x"67",x"71",x"E7",x"A4",x"22",x"3A",x"7A",x"64",x"47",x"03",x"70",x"77",x"5F",x"A1",x"DE",x"0F",x"58",x"10",x"50",x"06",x"FE",x"0C",x"6D",x"D7",x"89",x"E3",x"1C",x"64",x"50",x"A2",x"73",x"3A",x"0C",x"20",x"00",x"94",x"40",x"13",x"D5",x"C9",x"77",x"08",x"68",x"B8",x"6F",x"75",x"F3",x"0D",x"2C",x"58",x"18",x"44",x"61",x"73",x"0F",x"59",x"DC",x"63",x"B1",x"74",x"72",x"79",x"1B",x"AA",x"10",x"1D",x"E0",x"29",x"A1",x"34",x"72",x"65",x"3E",x"9B",x"42",x"42",x"74",x"A5",x"73",x"0F",x"62",x"6F",x"B5",x"72",x"D2",x"69",x"6E",x"D7",x"67",x"10",x"19",x"9F",x"86",x"76",x"4E",x"D1",x"CC",x"58",x"4D",x"66",x"75",x"A7",x"6C",x"97",x"73",x"8E",x"A8",x"64",x"20",x"FD",x"78",x"69",x"74",x"00",x"7A",x"1E",x"06",x"A2",x"61",x"6E",x"63",x"E8",x"65",x"6C",x"D3",x"00",x"8C",x"91",x"83",x"FB",x"B6",x"0B",x"11",x"06",x"10",x"40",x"10",x"02",x"6F",x"6B",x"FC",x"12",x"11",x"D1",x"47",x"E0",x"87",x"7C",x"A3",x"8A",x"FA",x"18",x"D0",x"78",x"20",x"89",x"FB",x"31",x"10",x"6B",x"F7",x"71",x"AD",x"F8",x"75",x"FD",x"68",x"F9",x"2D",x"0D",x"2F",x"FA",x"FB",x"B6",x"AD",x"29",x"64",x"7A",x"40",x"DF",x"AD",x"F8",x"02",x"90",x"05",x"DC",x"9F",x"55",x"CC",x"B6",x"12",x"DC",x"35",x"E3",x"40",x"B8",x"49",x"68",x"CE",x"15",x"FD",x"03",x"33",x"B6",x"16",x"47",x"14",x"5A",x"CD",x"D0",x"04",x"98",x"97",x"42",x"47",x"78",x"0A",x"79",x"9C",x"56",x"BC",x"33",x"38",x"3F",x"68",x"13",x"16",x"2C",x"BB",x"6C",x"8C",x"3F",x"58",x"78",x"58",x"47",x"F0",x"1A",x"E1",x"A1",x"1A",x"53",x"ED",x"12",x"1A",x"01",x"E5",x"1F",x"52",x"29",x"F0",x"1A",x"DA",x"AD",x"56",x"35",x"DF",x"83",x"57",x"48",x"A9",x"01",x"3A",x"09",x"46",x"A3",x"53",x"E6",x"7A",x"22",x"6D",x"1F",x"32",x"D6",x"28",x"05",x"23",x"E6",x"9D",x"DE",x"D0",x"BA",x"C4",x"7E",x"9D",x"E6",x"C9",x"F8",x"D0",x"EF",x"0E",x"53",x"0B",x"13",x"0E",x"DF",x"09",x"0A",x"91",x"A1",x"9A",x"85",x"91",x"71",x"DB",x"9F",x"DE",x"1D",x"3B",x"F3",x"60",x"67",x"62",x"9D",x"14",x"B4",x"F1",x"E5",x"6F",x"3C",x"F4",x"7C",x"CE",x"C2",x"F2",x"48",x"8F",x"96",x"24",x"13",x"F7",x"39",x"A2",x"5F",x"05",x"05",x"22",x"1F",x"A8",x"1D",x"A3",x"C6",x"C9",x"C4",x"DA",x"D3",x"13",x"A9",x"25",x"BD",x"A5",x"A4",x"48",x"4D",x"2B",x"D0",x"B5",x"8E",x"EC",x"A3",x"97",x"9E",x"A7",x"F0",x"1D",x"ED",x"19",x"ED",x"23",x"D2",x"E2",x"C7",x"39",x"2D",x"E5",x"44",x"2D",x"06",x"27",x"D4",x"A8",x"20",x"E6",x"1F",x"4C",x"9F",x"11",x"20",x"A8",x"FE",x"12",x"4F",x"EB",x"FB",x"95",x"AA",x"49",x"F6",x"EE",x"57",x"F3",x"78",x"DF",x"24",x"4F",x"8A",x"50",x"AA",x"54",x"F3",x"51",x"A7",x"0D",x"4F",x"2C",x"D0",x"49",x"11",x"04",x"A2",x"A6",x"86",x"08",x"58",x"C1",x"77",x"48",x"88",x"B5",x"EB",x"05",x"CA",x"00",x"24",x"A4",x"01",x"BE",x"1B",x"9E",x"AE",x"4E",x"BD",x"08",x"FF",x"AC",x"87",x"4C",x"0A",x"13",x"DA",x"9C",x"43",x"74",x"60",x"AE",x"9F",x"05",x"70",x"5D",x"F1",x"8E",x"58",x"E2",x"8A",x"A4",x"C0",x"CF",x"58",x"30",x"59",x"DE",x"31",x"7B",x"5A",x"32",x"EF",x"5B",x"33",x"BD",x"5C",x"F7",x"34",x"5D",x"DE",x"BD",x"35",x"E9",x"61",x"5E",x"45",x"5A",x"75",x"A5",x"AC",x"59",x"08",x"CE",x"21",x"D0",x"D3",x"0D",x"C2",x"78",x"C3",x"54",x"5A",x"80",x"AC",x"01",x"6C",x"EF",x"C0",x"8E",x"3D",x"B9",x"ED",x"99",x"B4",x"97",x"88",x"96",x"2C",x"F4",x"22",x"D2",x"6A",x"DE",x"4E",x"EF",x"04",x"2D",x"20",x"79",x"C6",x"13",x"02",x"AB",x"41",x"6C",x"A5",x"42",x"4E",x"EA",x"A9",x"81",x"27",x"F4",x"04",x"F2",x"C1",x"11",x"95",x"12",x"47",x"7A",x"C3",x"DE",x"0A",x"BD",x"C9",x"DF",x"FA",x"E8",x"93",x"D0",x"F1",x"91",x"BB",x"1F",x"5F",x"AD",x"84",x"0D",x"97",x"CA",x"B6",x"7B",x"5A",x"AA",x"55",x"58",x"6D",x"49",x"C1",x"55",x"F7",x"B6",x"AA",x"00",x"94",x"72",x"5E",x"73",x"A2",x"5B",x"DA",x"DE",x"E5",x"FA",x"52",x"64",x"7F",x"66",x"C7",x"B4",x"82",x"F4",x"4C",x"2E",x"44",x"06",x"C0",x"F3",x"CB",x"CD",x"03",x"3F",x"20",x"2C",x"14",x"12",x"BF",x"07",x"B5",x"08",x"F2",x"BB",x"AA",x"B5",x"08",x"F1",x"BB",x"2C",x"B6",x"DC",x"32",x"A2",x"F0",x"AB",x"6A",x"8B",x"B0",x"F3",x"AB",x"72",x"8B",x"B0",x"F4",x"AB",x"7A",x"8B",x"C1",x"B0",x"8D",x"F5",x"C3",x"7F",x"6E",x"14",x"E5",x"1D",x"57",x"A0",x"93",x"A3",x"18",x"32",x"99",x"63",x"A8",x"64",x"D0",x"BD",x"04",x"5B",x"17",x"5C",x"2C",x"0C",x"1B",x"39",x"C8",x"99",x"38",x"03",x"4D",x"D7",x"D0",x"C0",x"91",x"5E",x"A4",x"FD",x"BC",x"CA",x"D0",x"F8",x"9F",x"64",x"78",x"F2",x"E8",x"01",x"E5",x"2A",x"C8",x"F5",x"0A",x"4A",x"27",x"76",x"05",x"CD",x"C6",x"F0",x"26",x"DB",x"C7",x"C5",x"04",x"C8",x"13",x"C9",x"24",x"50",x"84",x"8D",x"9D",x"CA",x"45",x"4C",x"CB",x"80",x"A5",x"C8",x"AD",x"C7",x"1F",x"60",x"15",x"5C",x"92",x"B0",x"2C",x"59",x"46",x"62",x"63",x"F8",x"75",x"E5",x"5B",x"68",x"10",x"1C",x"1B",x"6D",x"D6",x"14",x"EB",x"37",x"A3",x"D7",x"B9",x"3E",x"59",x"C7",x"58",x"E3",x"04",x"F1",x"5A",x"78",x"59",x"34",x"32",x"58",x"C2",x"AD",x"B6",x"E9",x"35",x"56",x"DB",x"74",x"4D",x"55",x"9B",x"EA",x"CA",x"5A",x"9D",x"20",x"7A",x"5B",x"21",x"EF",x"5C",x"9D",x"73",x"CA",x"8D",x"5D",x"0D",x"E7",x"FC",x"A2",x"95",x"6C",x"EA",x"4D",x"DE",x"D6",x"88",x"F3",x"FA",x"AB",x"4A",x"6A",x"67",x"F5",x"AB",x"5A",x"12",x"B7",x"9F",x"60",x"B6",x"45",x"82",x"49",x"AA",x"DD",x"31",x"AD",x"92",x"C5",x"B2",x"AB",x"06",x"A1",x"27",x"4C",x"9C",x"C2",x"15",x"A5",x"BF",x"F7",x"8C",x"D6",x"60",x"AD",x"5E",x"A4",x"BE",x"AA",x"07",x"9C",x"E5",x"CD",x"00",x"DF",x"C0",x"0B",x"5E",x"53",x"4D",x"A2",x"27",x"BD",x"5D",x"0A",x"60",x"FD",x"7B",x"9D",x"C0",x"07",x"CA",x"BC",x"F2",x"D0",x"FE",x"8A",x"8F",x"FE",x"F0",x"06",x"F7",x"42",x"4C",x"EF",x"15",x"5E",x"DF",x"A6",x"CC",x"3E",x"53",x"1F",x"38",x"6B",x"50",x"DE",x"07",x"EE",x"56",x"5E",x"B4",x"29",x"2A",x"EF",x"01",x"7C",x"52",x"DE",x"03",x"F8",x"88",x"F2",x"1E",x"C0",x"27",x"E5",x"15",x"01",x"BA",x"94",x"CA",x"CB",x"00",x"CE",x"A5",x"F2",x"BC",x"4A",x"54",x"0A",x"37",x"60",x"79",x"1B",x"68",x"6F",x"24",x"FC",x"0E",x"AF",x"A9",x"0E",x"CB",x"BF",x"9D",x"A9",x"21",x"2F",x"CD",x"A2",x"AC",x"DA",x"86",x"DF",x"03",x"B0",x"1D",x"00",x"BF",x"0C",x"16",x"69",x"C8",x"04",x"12",x"BF",x"39",x"32",x"31",x"98",x"5A",x"2C",x"3F",x"F4",x"FB",x"40",x"59",x"33",x"5B",x"31",x"91",x"47",x"9B",x"EB",x"63",x"7F",x"0D",x"18",x"09",x"E7",x"A5",x"4D",x"19",x"6D",x"2B",x"37",x"CC",x"C8",x"60",x"7D",x"D2",x"0C",x"74",x"98",x"18",x"6D",x"FC",x"D6",x"A8",x"F6",x"C2",x"10",x"66",x"98",x"49",x"9A",x"09",x"94",x"66",x"8D",x"0A",x"16",x"FB",x"2B",x"68",x"0A",x"2A",x"A4",x"75",x"70",x"09",x"C0",x"D2",x"40",x"18",x"60",x"DD",x"A6",x"C2",x"AD",x"A9",x"C2",x"F9",x"BE",x"0B",x"64",x"23",x"0A",x"BB",x"A5",x"94",x"AE",x"13",x"60",x"EE",x"5E",x"AD",x"B2",x"64",x"F0",x"F8",x"33",x"34",x"10",x"D6",x"D3",x"28",x"82",x"14",x"4E",x"94",x"82",x"4F",x"0E",x"72",x"D0",x"59",x"98",x"CA",x"18",x"E7",x"E0",x"C3",x"05",x"4A",x"4B",x"8B",x"66",x"87",x"3E",x"1A",x"DC",x"28",x"F9",x"DD",x"0F",x"E4",x"47",x"C2",x"AE",x"A1",x"74",x"C1",x"75",x"E2",x"28",x"E1",x"02",x"91",x"6E",x"E6",x"E9",x"23",x"8A",x"B3",x"1D",x"70",x"8F",x"29",x"1D",x"C1",x"90",x"10",x"85",x"FC",x"F3",x"D6",x"E2",x"09",x"AE",x"08",x"F6",x"83",x"D7",x"55",x"E3",x"39",x"F7",x"DD",x"61",x"47",x"3D",x"8F",x"F7",x"08",x"20",x"E4",x"71",x"B0",x"51",x"4C",x"D2",x"D5",x"A0",x"5F",x"12",x"8C",x"CF",x"1B",x"C2",x"10",x"8F",x"C8",x"05",x"89",x"30",x"48",x"AD",x"01",x"71",x"FB",x"A8",x"F7",x"B6",x"8C",x"4A",x"6A",x"9B",x"DF",x"00",x"2F",x"90",x"A5",x"C6",x"68",x"A8",x"64",x"B1",x"A4",x"FF",x"4D",x"65",x"99",x"2D",x"15",x"76",x"15",x"DB",x"CA",x"E3",x"62",x"17",x"84",x"0D",x"2C",x"4C",x"35",x"DC",x"19",x"AD",x"E3",x"D5",x"CD",x"BC",x"A0",x"0A",x"20",x"D5",x"04",x"43",x"26",x"55",x"30",x"B2",x"32",x"A2",x"89",x"D9",x"5A",x"77",x"C8",x"D6",x"CD",x"00",x"E1",x"EC",x"06",x"C4",x"52",x"EA",x"05",x"37",x"26",x"D0",x"8B",x"9D",x"18",x"4C",x"63",x"E7",x"EF",x"AB",x"C0",x"AD",x"0B",x"5A",x"3A",x"1E",x"03",x"30",x"B0",x"11",x"F8",x"A6",x"54",x"20",x"B8",x"D1",x"17",x"8C",x"9F",x"E3",x"D1",x"91",x"50",x"E6",x"77",x"B1",x"93",x"FB",x"59",x"30",x"AC",x"5B",x"91",x"A5",x"9D",x"F3",x"F6",x"EE",x"BF",x"05",x"53",x"4F",x"A3",x"3B",x"E8",x"AC",x"07",x"16",x"18",x"71",x"1F",x"7C",x"05",x"6A",x"45",x"02",x"AD",x"46",x"75",x"2C",x"58",x"DC",x"02",x"48",x"CF",x"ED",x"5C",x"41",x"3E",x"AC",x"0B",x"B8",x"66",x"3C",x"08",x"6E",x"14",x"C5",x"98",x"1A",x"16",x"07",x"1C",x"99",x"CE",x"90",x"1D",x"C5",x"50",x"63",x"1F",x"07",x"68",x"9D",x"A9",x"B0",x"AD",x"6F",x"71",x"9A",x"6D",x"1D",x"BE",x"6C",x"D9",x"D6",x"FD",x"1A",x"60",x"DB",x"2A",x"42",x"1B",x"A6",x"B2",x"F0",x"E0",x"96",x"E7",x"61",x"A9",x"92",x"6D",x"7B",x"B5",x"0E",x"81",x"56",x"D6",x"07",x"24",x"6D",x"35",x"7C",x"C0",x"1B",x"DE",x"F3",x"20",x"6D",x"CF",x"99",x"42",x"43",x"32",x"97",x"2C",x"A4",x"ED",x"B9",x"ED",x"46",x"2F",x"C5",x"F8",x"B7",x"C7",x"2C",x"A3",x"81",x"4F",x"A0",x"C7",x"D9",x"FF",x"60",x"3C",x"F2",x"D7",x"91",x"13",x"60",x"A0",x"09",x"17",x"EE",x"CC",x"F8",x"54",x"06",x"E5",x"97",x"2C",x"BC",x"5A",x"F4",x"65",x"D9",x"10",x"D9",x"1A",x"E0",x"0D",x"A0",x"5E",x"F0",x"18",x"AE",x"0D",x"1A",x"8D",x"D8",x"63",x"33",x"A3",x"B9",x"47",x"46",x"20",x"C1",x"04",x"07",x"2B",x"06",x"90",x"BF",x"0B",x"10",x"4C",x"C2",x"4A",x"C6",x"A0",x"61",x"17",x"F0",x"D1",x"11",x"38",x"57",x"05",x"58",x"02",x"B6",x"6F",x"1D",x"C2",x"20",x"89",x"2D",x"B0",x"F2",x"36",x"56",x"EF",x"85",x"B4",x"A0",x"F9",x"08",x"73",x"86",x"3C",x"4D",x"FE",x"36",x"9A",x"40",x"DD",x"3F",x"6C",x"13",x"79",x"55",x"02",x"16",x"1B",x"64",x"E4",x"C1",x"23",x"1F",x"9C",x"95",x"24",x"8E",x"39",x"72",x"1A",x"D9",x"50",x"92",x"DC",x"32",x"E2",x"40",x"36",x"3A",x"01",x"AE",x"45",x"7E",x"09",x"BD",x"0A",x"75",x"CB",x"5A",x"9D",x"21",x"19",x"0F",x"D9",x"08",x"BA",x"08",x"48",x"1D",x"D7",x"55",x"0C",x"EA",x"05",x"93",x"D6",x"3C",x"4C",x"9A",x"F7",x"1C",x"31",x"42",x"4F",x"B0",x"2D",x"DF",x"AA",x"CA",x"0A",x"B6",x"65",x"B3",x"AA",x"0E",x"DD",x"B7",x"01",x"1C",x"90",x"02",x"80",x"18",x"7F",x"73",x"14",x"E5",x"10",x"6C",x"12",x"5A",x"68",x"06",x"39",x"48",x"C9",x"34",x"B0",x"04",x"68",x"FD",x"88",x"DF",x"1C",x"4F",x"B2",x"AA",x"5E",x"D1",x"33",x"C7",x"8A",x"86",x"4E",x"8D",x"53",x"76",x"21",x"A4",x"D2",x"3A",x"60",x"C1",x"E1",x"99",x"DB",x"62",x"AF",x"6C",x"29",x"A8",x"9F",x"D0",x"65",x"35",x"1C",x"C9",x"DA",x"61",x"0E",x"36",x"A4",x"B2",x"61",x"98",x"0B",x"44",x"D3",x"9D",x"6D",x"1C",x"55",x"DF",x"C0",x"02",x"57",x"DB",x"20",x"21",x"1D",x"80",x"D6",x"FD",x"14",x"73",x"DC",x"90",x"B7",x"87",x"00",x"1F",x"1C",x"09",x"49",x"12",x"A0",x"44",x"5E",x"E0",x"60",x"B2",x"7D",x"4D",x"C0",x"A3",x"82",x"D1",x"28",x"02",x"2A",x"83",x"51",x"38",x"58",x"1C",x"69",x"8D",x"4D",x"06",x"5F",x"45",x"0F",x"89",x"04",x"45",x"85",x"80",x"0D",x"E0",x"03",x"40",x"22",x"1B",x"40",x"53",x"50",x"80",x"9B",x"64",x"49",x"12",x"45",x"C2",x"74",x"F9",x"39",x"6F",x"9D",x"CE",x"CF",x"1D",x"A7",x"09",x"40",x"F1",x"21",x"A0",x"02",x"2C",x"B8",x"02",x"81",x"43",x"1B",x"88",x"98",x"44",x"80",x"89",x"18",x"08",x"B2",x"56",x"29",x"BF",x"EA",x"E9",x"92",x"F7",x"20",x"6F",x"1D",x"A3",x"7F",x"07",x"28",x"7E",x"40",x"56",x"4F",x"C2",x"BD",x"72",x"D5",x"04",x"89",x"4A",x"75",x"3B",x"CA",x"29",x"1E",x"AA",x"79",x"30",x"1A",x"AD",x"3A",x"75",x"0F",x"D2",x"E8",x"F8",x"12",x"C9",x"67",x"B0",x"0E",x"FC",x"37",x"6B",x"48",x"E9",x"30",x"D9",x"20",x"CD",x"1E",x"F8",x"F7",x"23",x"22",x"05",x"5A",x"20",x"E0",x"9A",x"15",x"7A",x"99",x"BF",x"7B",x"9D",x"33",x"4C",x"9F",x"3C",x"1E",x"97",x"E5",x"C9",x"68",x"65",x"41",x"03",x"5C",x"28",x"A4",x"09",x"02",x"A5",x"38",x"2E",x"AA",x"E9",x"A5",x"D6",x"2F",x"53",x"99",x"0D",x"60",x"C7",x"96",x"EA",x"69",x"75",x"49",x"13",x"96",x"87",x"7B",x"F0",x"13",x"25",x"3E",x"30",x"01",x"B9",x"8F",x"1A",x"20",x"67",x"84",x"16",x"93",x"FC",x"44",x"41",x"0F",x"88",x"0C",x"C6",x"95",x"8E",x"B3",x"58",x"70",x"6A",x"02",x"60",x"E9",x"11",x"1F",x"41",x"57",x"A4",x"17",x"8C",x"71",x"8A",x"CE",x"96",x"2E",x"00",x"B3",x"F0",x"DD",x"06",x"47",x"EE",x"45",x"4C",x"ED",x"1E",x"20",x"36",x"1F",x"FF",x"D9",x"38",x"F0",x"86",x"13",x"37",x"26",x"B3",x"A5",x"CE",x"B2",x"C9",x"06",x"F0",x"08",x"BF",x"02",x"1E",x"4C",x"16",x"1F",x"F2",x"B1",x"A6",x"68",x"89",x"50",x"82",x"05",x"35",x"61",x"5A",x"C0",x"8C",x"AD",x"48",x"76",x"4A",x"8D",x"A2",x"59",x"25",x"83",x"4A",x"78",x"3F",x"2F",x"DB",x"C5",x"E6",x"B3",x"18",x"1D",x"D5",x"65",x"34",x"B4",x"96",x"40",x"14",x"52",x"B6",x"AF",x"CA",x"68",x"D4",x"54",x"4E",x"7C",x"80",x"B0",x"FE",x"78",x"77",x"1F",x"5F",x"E4",x"AD",x"E5",x"31",x"5A",x"35",x"CE",x"74",x"65",x"3E",x"04",x"47",x"E6",x"B8",x"AC",x"A5",x"8D",x"26",x"A7",x"C5",x"61",x"0B",x"A3",x"C9",x"69",x"CD",x"D8",x"C2",x"CA",x"A6",x"F8",x"F0",x"32",x"83",x"BA",x"3A",x"8E",x"9D",x"21",x"C6",x"AC",x"B1",x"B4",x"11",x"22",x"AA",x"51",x"23",x"CA",x"D4",x"2D",x"A6",x"D1",x"54",x"E9",x"3D",x"A5",x"15",x"E9",x"9E",x"B5",x"C7",x"AA",x"A9",x"A0",x"E8",x"91",x"A8",x"6B",x"28",x"A7",x"B1",x"B0",x"52",x"E7",x"60",x"30",x"0B",x"6B",x"0F",x"DA",x"25",x"94",x"A9",x"0A",x"1C",x"F1",x"0F",x"0F",x"49",x"2C",x"18",x"69",x"01",x"3A",x"40",x"0A",x"A1",x"D2",x"42",x"8E",x"15",x"4C",x"4C",x"D8",x"4A",x"0B",x"AD",x"4D",x"96",x"FF",x"7D",x"39",x"0D",x"58",x"50",x"8D",x"11",x"4E",x"9D",x"00",x"F0",x"21",x"E9",x"76",x"8B",x"51",x"03",x"53",x"D6",x"CA",x"CB",x"FF",x"5E",x"D9",x"A5",x"47",x"4E",x"76",x"00",x"F5",x"90",x"8C",x"A0",x"D1",x"92",x"AF",x"6E",x"62",x"42",x"B5",x"43",x"46",x"01",x"B3",x"EB",x"A6",x"1F",x"6D",x"E0",x"90",x"0E",x"AE",x"BA",x"EC",x"B0",x"12",x"D0",x"F0",x"FB",x"36",x"1F",x"5E",x"4C",x"36",x"EE",x"AD",x"C7",x"B5",x"2E",x"0A",x"2E",x"07",x"7E",x"2B",x"40",x"D6",x"EA",x"EA",x"3A",x"4C",x"20",x"BC",x"0C",x"AF",x"C8",x"80",x"C9",x"F7",x"CA",x"8A",x"CB",x"EA",x"2A",x"72",x"41",x"79",x"53",x"42",x"AD",x"8D",x"CF",x"D6",x"4C",x"BE",x"FF",x"6E",x"05",x"05",x"97",x"36",x"42",x"A4",x"07",x"15",x"F4",x"13",x"9D",x"0B",x"16",x"3A",x"9A",x"A5",x"08",x"EC",x"AD",x"8A",x"BE",x"00",x"0A",x"97",x"D8",x"55",x"20",x"C7",x"17",x"D4",x"F4",x"5B",x"08",x"FF",x"BB",x"85",x"46",x"1F",x"67",x"1E",x"91",x"1E",x"BB",x"1E",x"E5",x"1E",x"0F",x"56",x"19",x"39",x"0E",x"63",x"AB",x"7F",x"53",x"63",x"00",x"39",x"78",x"01",x"E7",x"A2",x"02",x"9C",x"CC",x"F3",x"20",x"03",x"97",x"F6",x"21",x"5C",x"16",x"3A",x"04",x"55",x"2B",x"C6",x"9F",x"F1",x"4A",x"22",x"0D",x"6A",x"4E",x"70",x"0E",x"26",x"31",x"E0",x"3A",x"06",x"8C",x"4A",x"C0",x"24",x"04",x"06",x"3C",x"0E",x"1C",x"07",x"DC",x"81",x"0F",x"33",x"03",x"0E",x"0F",x"14",x"13",x"02",x"74",x"9C",x"09",x"14",x"78",x"1A",x"18",x"8F",x"81",x"10",x"33",x"03",x"1A",x"0F",x"21",x"23",x"0C",x"30",x"69",x"A2",x"01",x"4F",x"18",x"6E",x"A0",x"24",x"B0",x"8C",x"6E",x"81",x"C0",x"28",x"D0",x"E7",x"F9",x"63",x"4C",x"48",x"01",x"AD",x"49",x"B5",x"20",x"8E",x"B0",x"A9",x"11",x"85",x"B1",x"7B",x"7E",x"7D",x"78",x"A8",x"65",x"D5",x"67",x"7C",x"AC",x"9B",x"CD",x"B5",x"D0",x"6C",x"98",x"88",x"51",x"18",x"78",x"75",x"71",x"79",x"A8",x"06",x"3A",x"CD",x"A0",x"F0",x"B0",x"54",x"D7",x"A2",x"07",x"28",x"91",x"3F",x"A5",x"21",x"2F",x"C6",x"DB",x"1B",x"23",x"0A",x"E3",x"30",x"15",x"26",x"E7",x"8C",x"0D",x"3C",x"F2",x"0E",x"60",x"81",x"83",x"54",x"60",x"40",x"7F",x"1F",x"4A",x"51",x"11",x"3D",x"12",x"12",x"39",x"76",x"C0",x"13",x"3B",x"26",x"14",x"93",x"32",x"0B",x"A2",x"02",x"4A",x"39",x"EA",x"0C",x"6A",x"91",x"51",x"75",x"A9",x"D3",x"AE",x"EF",x"6D",x"81",x"8D",x"92",x"20",x"58",x"23",x"EC",x"77",x"D7",x"DD",x"04",x"B0",x"73",x"ED",x"0B",x"B5",x"56",x"F1",x"23",x"DC",x"F3",x"19",x"90",x"46",x"20",x"3D",x"24",x"87",x"1D",x"BA",x"1E",x"DF",x"8F",x"8D",x"64",x"CB",x"25",x"1D",x"49",x"43",x"6E",x"1D",x"E7",x"19",x"15",x"9C",x"08",x"11",x"A8",x"CD",x"CA",x"E3",x"39",x"D0",x"F8",x"2E",x"98",x"D6",x"2D",x"67",x"8A",x"48",x"47",x"53",x"F7",x"F0",x"8B",x"E7",x"E2",x"01",x"6D",x"06",x"0C",x"41",x"AA",x"B7",x"23",x"51",x"83",x"F0",x"D0",x"25",x"AD",x"74",x"F8",x"22",x"38",x"ED",x"0E",x"C9",x"21",x"A8",x"4C",x"4F",x"4C",x"EB",x"23",x"EA",x"A9",x"10",x"2F",x"20",x"BC",x"ED",x"26",x"AF",x"19",x"08",x"00",x"67",x"0F",x"71",x"01",x"16",x"15",x"02",x"67",x"1B",x"71",x"03",x"12",x"22",x"B0",x"62",x"56",x"04",x"25",x"C9",x"24",x"90",x"17",x"A9",x"EA",x"05",x"4C",x"2B",x"24",x"60",x"C5",x"FF",x"F0",x"95",x"D0",x"BF",x"2C",x"21",x"53",x"AD",x"76",x"22",x"F0",x"25",x"5A",x"0C",x"7C",x"EB",x"C2",x"C9",x"A0",x"4F",x"EB",x"2F",x"8F",x"24",x"B5",x"5C",x"F3",x"F0",x"20",x"55",x"27",x"AE",x"44",x"A8",x"06",x"15",x"1A",x"C8",x"70",x"A0",x"58",x"86",x"3A",x"85",x"FA",x"20",x"96",x"31",x"BF",x"F0",x"49",x"90",x"9D",x"94",x"18",x"45",x"E0",x"05",x"F1",x"4A",x"46",x"4A",x"19",x"03",x"B5",x"49",x"CA",x"D3",x"86",x"48",x"17",x"33",x"66",x"21",x"E8",x"A3",x"E8",x"D0",x"ED",x"00",x"4D",x"E0",x"80",x"57",x"08",x"44",x"E0",x"CB",x"D6",x"6F",x"5A",x"AA",x"47",x"02",x"D3",x"CA",x"B6",x"02",x"A2",x"13",x"9E",x"10",x"E0",x"0C",x"EC",x"8A",x"AB",x"4B",x"04",x"9E",x"D2",x"E2",x"DF",x"25",x"1F",x"11",x"B0",x"12",x"91",x"72",x"92",x"2C",x"0C",x"33",x"A7",x"94",x"5F",x"EB",x"E2",x"2E",x"37",x"EE",x"31",x"30",x"19",x"EB",x"11",x"09",x"9C",x"E9",x"74",x"71",x"52",x"07",x"B9",x"52",x"74",x"25",x"87",x"20",x"6D",x"26",x"DD",x"DE",x"00",x"E0",x"1C",x"C1",x"00",x"3D",x"A0",x"F0",x"B1",x"AA",x"75",x"B4",x"1D",x"64",x"00",x"88",x"73",x"57",x"C0",x"3E",x"78",x"1F",x"F0",x"8C",x"00",x"78",x"06",x"D8",x"6A",x"98",x"59",x"2E",x"4D",x"82",x"03",x"85",x"06",x"48",x"16",x"2B",x"34",x"58",x"B2",x"B4",x"B3",x"F5",x"C1",x"00",x"61",x"14",x"8B",x"A5",x"A7",x"D0",x"1F",x"87",x"B3",x"F0",x"01",x"67",x"89",x"95",x"5D",x"91",x"A8",x"60",x"B8",x"3E",x"0A",x"A3",x"9A",x"C9",x"24",x"03",x"16",x"DF",x"50",x"8A",x"BD",x"85",x"AD",x"B1",x"44",x"A8",x"2C",x"08",x"A2",x"A9",x"BA",x"F0",x"06",x"C8",x"E8",x"E4",x"AD",x"FC",x"D0",x"F6",x"86",x"8C",x"AF",x"38",x"FB",x"C4",x"1F",x"AA",x"22",x"2D",x"AB",x"38",x"C7",x"01",x"E5",x"BE",x"AD",x"27",x"AC",x"8D",x"D7",x"E2",x"A5",x"42",x"72",x"04",x"05",x"37",x"49",x"E8",x"A8",x"D4",x"37",x"01",x"14",x"4E",x"A7",x"BB",x"E9",x"A9",x"B3",x"E3",x"CE",x"68",x"48",x"11",x"DA",x"F9",x"03",x"20",x"90",x"47",x"B9",x"F7",x"B9",x"00",x"4A",x"C4",x"00",x"D4",x"5C",x"FE",x"8E",x"68",x"48",x"11",x"3D",x"91",x"FB",x"AA",x"34",x"9D",x"11",x"AA",x"18",x"D9",x"65",x"95",x"05",x"A9",x"58",x"1E",x"B5",x"3C",x"6E",x"FE",x"28",x"4C",x"B4",x"42",x"40",x"4C",x"27",x"8B",x"54",x"A9",x"A2",x"D1",x"48",x"8B",x"84",x"68",x"5D",x"28",x"3D",x"EA",x"60",x"ED",x"20",x"19",x"89",x"51",x"A7",x"72",x"53",x"30",x"BA",x"5E",x"21",x"A1",x"EB",x"1B",x"89",x"B1",x"28",x"14",x"36",x"D5",x"A0",x"FF",x"84",x"42",x"F3",x"53",x"0A",x"A8",x"B7",x"41",x"40",x"72",x"92",x"B0",x"48",x"F0",x"FA",x"36",x"C9",x"36",x"D4",x"A9",x"36",x"38",x"B7",x"0F",x"70",x"07",x"84",x"44",x"C2",x"6F",x"72",x"DF",x"5D",x"24",x"72",x"29",x"BB",x"90",x"03",x"4C",x"23",x"28",x"18",x"98",x"65",x"FF",x"39",x"A1",x"38",x"81",x"44",x"52",x"B9",x"16",x"D4",x"7B",x"4C",x"92",x"27",x"2A",x"F7",x"E0",x"14",x"E3",x"CD",x"01",x"AB",x"E8",x"4C",x"BE",x"27",x"F8",x"45",x"5A",x"05",x"47",x"16",x"99",x"BD",x"02",x"5A",x"06",x"5C",x"EB",x"09",x"01",x"BD",x"AB",x"3A",x"6A",x"2B",x"0A",x"0A",x"0A",x"D1",x"1E",x"AD",x"4E",x"3B",x"51",x"46",x"0F",x"02",x"2B",x"54",x"96",x"29",x"3E",x"01",x"85",x"47",x"EE",x"49",x"22",x"45",x"20",x"34",x"4B",x"12",x"AB",x"4C",x"17",x"28",x"43",x"A7",x"C7",x"E0",x"EF",x"E2",x"0B",x"86",x"C2",x"42",x"AD",x"5B",x"FF",x"2D",x"31",x"DC",x"13",x"A8",x"25",x"C7",x"0A",x"8D",x"6E",x"F5",x"10",x"1C",x"ED",x"0D",x"84",x"4C",x"3C",x"28",x"F6",x"27",x"3A",x"7A",x"A9",x"0C",x"FD",x"41",x"4F",x"D4",x"03",x"84",x"CE",x"43",x"8A",x"A8",x"27",x"F0",x"13",x"7B",x"B6",x"B1",x"EA",x"92",x"CE",x"ED",x"A4",x"43",x"CE",x"31",x"C8",x"4C",x"40",x"28",x"F9",x"D7",x"E8",x"F5",x"35",x"F4",x"13",x"60",x"A6",x"46",x"07",x"4A",x"98",x"04",x"A6",x"CE",x"0C",x"20",x"06",x"02",x"33",x"09",x"D0",x"ED",x"A0",x"49",x"B4",x"2A",x"6A",x"88",x"6D",x"82",x"B6",x"40",x"64",x"68",x"12",x"D3",x"F5",x"08",x"70",x"26",x"4C",x"F8",x"28",x"E0",x"06",x"D0",x"1D",x"FF",x"EB",x"3A",x"09",x"04",x"27",x"92",x"2C",x"3A",x"FB",x"A9",x"0A",x"21",x"7A",x"3C",x"20",x"F2",x"D2",x"2F",x"06",x"AB",x"A2",x"FF",x"60",x"E8",x"49",x"F5",x"30",x"E7",x"CE",x"A5",x"BA",x"9A",x"D8",x"31",x"BE",x"33",x"E5",x"07",x"60",x"1F",x"78",x"AD",x"14",x"43",x"FB",x"C5",x"5A",x"FC",x"C8",x"91",x"97",x"18",x"A9",x"02",x"65",x"3E",x"34",x"FD",x"A5",x"3D",x"FE",x"9A",x"84",x"DE",x"B3",x"E5",x"83",x"8B",x"76",x"B9",x"44",x"34",x"85",x"0F",x"30",x"D2",x"26",x"BD",x"29",x"53",x"40",x"C6",x"D6",x"E7",x"A9",x"B7",x"FF",x"91",x"86",x"50",x"BA",x"5C",x"2A",x"E4",x"B2",x"E9",x"2C",x"90",x"2B",x"49",x"7D",x"70",x"D0",x"04",x"47",x"FE",x"2D",x"49",x"ED",x"70",x"FB",x"93",x"39",x"B8",x"1A",x"C8",x"8A",x"48",x"C7",x"8A",x"8C",x"A0",x"21",x"29",x"14",x"48",x"49",x"01",x"7D",x"51",x"10",x"10",x"47",x"AA",x"C2",x"79",x"2F",x"D4",x"28",x"8E",x"17",x"8A",x"C3",x"45",x"6F",x"01",x"8F",x"8A",x"08",x"68",x"C8",x"CA",x"AA",x"E8",x"8E",x"7C",x"06",x"EC",x"ED",x"96",x"C2",x"BA",x"C2",x"21",x"07",x"10",x"95",x"0D",x"0B",x"F0",x"1F",x"98",x"95",x"04",x"18",x"26",x"02",x"60",x"A7",x"10",x"58",x"DD",x"30",x"8F",x"31",x"1A",x"6D",x"4E",x"A8",x"B5",x"09",x"16",x"B0",x"12",x"EE",x"00",x"16",x"71",x"D2",x"0F",x"AC",x"00",x"11",x"26",x"12",x"60",x"C7",x"3D",x"50",x"26",x"06",x"68",x"CD",x"C4",x"31",x"84",x"C5",x"52",x"A0",x"D7",x"48",x"67",x"0D",x"28",x"2B",x"E8",x"25",x"07",x"7A",x"93",x"26",x"62",x"04",x"49",x"30",x"D9",x"38",x"E9",x"D1",x"09",x"1F",x"1F",x"B0",x"09",x"EE",x"00",x"1F",x"A1",x"B2",x"02",x"A6",x"4C",x"0B",x"34",x"5E",x"E4",x"5F",x"15",x"89",x"60",x"AE",x"91",x"78",x"6B",x"D8",x"03",x"D3",x"53",x"6C",x"51",x"7C",x"85",x"1C",x"0B",x"A6",x"A0",x"15",x"60",x"D0",x"09",x"E4",x"B2",x"F0",x"0A",x"FF",x"5E",x"2A",x"30",x"05",x"BD",x"58",x"75",x"3D",x"E8",x"74",x"4B",x"2E",x"F5",x"F0",x"73",x"71",x"01",x"C0",x"08",x"BB",x"BC",x"3A",x"6F",x"CA",x"59",x"03",x"F8",x"C7",x"E7",x"49",x"81",x"D0",x"AC",x"EB",x"9A",x"47",x"EB",x"8B",x"11",x"60",x"64",x"8E",x"41",x"5A",x"E7",x"00",x"2C",x"2A",x"4B",x"41",x"E1",x"1D",x"18",x"97",x"4C",x"09",x"60",x"8E",x"E6",x"6D",x"E0",x"8E",x"3C",x"59",x"67",x"2D",x"C5",x"70",x"72",x"04",x"E8",x"75",x"AE",x"67",x"08",x"64",x"1F",x"63",x"12",x"66",x"65",x"62",x"02",x"FD",x"A3",x"56",x"01",x"D2",x"61",x"6C",x"07",x"6A",x"75",x"BF",x"06",x"74",x"72",x"03",x"D8",x"6D",x"61",x"79",x"05",x"6E",x"5F",x"76",x"11",x"6F",x"63",x"F4",x"74",x"10",x"73",x"65",x"70",x"BF",x"FF",x"04",x"03",x"07",x"F5",x"08",x"AA",x"06",x"05",x"01",x"0B",x"0A",x"09",x"02",x"76",x"7F",x"16",x"AE",x"1E",x"51",x"C2",x"08",x"1F",x"20",x"FF",x"E4",x"D3",x"8B",x"30",x"02",x"30",x"31",x"19",x"67",x"5C",x"E9",x"BC",x"A9",x"BF",x"99",x"69",x"80",x"13",x"32",x"41",x"0F",x"04",x"79",x"90",x"0A",x"13",x"34",x"FC",x"0E",x"24",x"F2",x"6E",x"73",x"C9",x"02",x"CB",x"35",x"AE",x"D2",x"F0",x"05",x"A2",x"01",x"F2",x"29",x"44",x"10",x"8E",x"22",x"A7",x"BD",x"29",x"03",x"F0",x"0D",x"F1",x"08",x"1D",x"11",x"4B",x"28",x"FE",x"8C",x"A0",x"C9",x"1E",x"90",x"F8",x"A9",x"FB",x"29",x"65",x"44",x"09",x"25",x"C6",x"53",x"22",x"2D",x"46",x"4D",x"63",x"BD",x"21",x"26",x"0E",x"AA",x"82",x"46",x"C9",x"0D",x"90",x"E2",x"05",x"99",x"12",x"3A",x"89",x"10",x"7E",x"43",x"01",x"CB",x"A1",x"1C",x"7D",x"D6",x"76",x"D6",x"92",x"ED",x"88",x"CD",x"53",x"65",x"90",x"0C",x"AE",x"EF",x"FF",x"EE",x"4D",x"8C",x"2C",x"24",x"56",x"60",x"A4",x"7A",x"D3",x"DF",x"93",x"8A",x"CC",x"6A",x"29",x"41",x"F0",x"16",x"C9",x"A0",x"B0",x"10",x"3F",x"40",x"4A",x"AA",x"F2",x"16",x"EF",x"5C",x"8F",x"AA",x"80",x"CC",x"02",x"A2",x"5A",x"AD",x"6F",x"C9",x"0A",x"B0",x"07",x"F6",x"8A",x"18",x"6D",x"27",x"AA",x"60",x"5B",x"09",x"69",x"25",x"FD",x"F2",x"BA",x"A2",x"20",x"69",x"9D",x"29",x"7A",x"37",x"FA",x"A6",x"DF",x"B4",x"9D",x"1B",x"42",x"93",x"AB",x"B3",x"E0",x"F0",x"0E",x"D1",x"37",x"AA",x"EB",x"13",x"24",x"7D",x"3B",x"D0",x"F5",x"A4",x"B3",x"FB",x"AD",x"03",x"99",x"B6",x"97",x"A3",x"A2",x"AD",x"21",x"C5",x"00",x"D5",x"45",x"DA",x"12",x"D9",x"79",x"2C",x"E5",x"F0",x"02",x"80",x"0B",x"87",x"6F",x"07",x"36",x"C8",x"C0",x"D4",x"33",x"EB",x"FA",x"6F",x"40",x"E8",x"88",x"C4",x"B3",x"D0",x"0E",x"FE",x"0A",x"F0",x"A5",x"CA",x"52",x"46",x"46",x"5E",x"99",x"FE",x"0C",x"1B",x"C2",x"0C",x"D0",x"F7",x"C6",x"38",x"87",x"6E",x"3D",x"72",x"20",x"26",x"2F",x"EF",x"F4",x"64",x"20",x"70",x"A2",x"0C",x"27",x"1D",x"64",x"7A",x"AC",x"5E",x"38",x"A3",x"2E",x"CA",x"D0",x"FA",x"47",x"E6",x"90",x"4D",x"06",x"1C",x"55",x"7B",x"A0",x"69",x"48",x"9B",x"DD",x"D8",x"E4",x"5B",x"28",x"E2",x"81",x"56",x"EA",x"11",x"B0",x"95",x"C0",x"5C",x"E1",x"BA",x"A1",x"20",x"51",x"2D",x"7A",x"6C",x"75",x"81",x"2F",x"FC",x"C8",x"5A",x"56",x"A3",x"92",x"F2",x"7F",x"3C",x"2C",x"2F",x"04",x"1B",x"E8",x"C2",x"03",x"D0",x"EF",x"BF",x"2D",x"53",x"A0",x"0E",x"3F",x"A5",x"C2",x"A7",x"E4",x"00",x"8C",x"67",x"7A",x"B6",x"54",x"4A",x"D0",x"05",x"60",x"FB",x"0D",x"91",x"0E",x"69",x"8D",x"B5",x"55",x"20",x"FD",x"2A",x"AC",x"F7",x"65",x"22",x"95",x"18",x"23",x"2A",x"3D",x"D1",x"74",x"C8",x"A6",x"AB",x"A5",x"44",x"09",x"70",x"9D",x"B1",x"BE",x"E6",x"43",x"68",x"EF",x"D5",x"03",x"A8",x"6E",x"B3",x"B1",x"98",x"21",x"B9",x"06",x"E2",x"35",x"50",x"AB",x"11",x"14",x"00",x"8A",x"43",x"2F",x"6D",x"1D",x"E8",x"29",x"AD",x"5C",x"08",x"B8",x"55",x"91",x"2B",x"65",x"6C",x"7E",x"D1",x"B2",x"83",x"CB",x"B2",x"0A",x"C9",x"23",x"DE",x"A0",x"4C",x"C4",x"E2",x"A9",x"AE",x"D1",x"EF",x"06",x"5A",x"98",x"AA",x"B2",x"8E",x"B3",x"B1",x"89",x"C8",x"AA",x"CA",x"BD",x"9C",x"8D",x"61",x"59",x"CC",x"AC",x"96",x"AD",x"21",x"2D",x"01",x"EE",x"20",x"DD",x"2F",x"6D",x"C8",x"1C",x"F6",x"E3",x"60",x"98",x"EF",x"48",x"45",x"65",x"87",x"B9",x"9A",x"7E",x"A6",x"AF",x"45",x"45",x"CB",x"8B",x"4A",x"44",x"F5",x"F7",x"46",x"01",x"A3",x"C5",x"DE",x"6B",x"04",x"FC",x"93",x"38",x"A9",x"28",x"E5",x"FF",x"4A",x"18",x"65",x"7A",x"E8",x"A4",x"04",x"A4",x"44",x"AF",x"64",x"BD",x"00",x"47",x"48",x"F4",x"89",x"DE",x"60",x"B6",x"88",x"A0",x"F1",x"04",x"90",x"84",x"0A",x"94",x"42",x"E8",x"03",x"23",x"56",x"F8",x"01",x"0C",x"4A",x"AD",x"5A",x"8D",x"68",x"4B",x"57",x"15",x"39",x"18",x"93",x"80",x"02",x"4A",x"51",x"04",x"30",x"BD",x"01",x"55",x"46",x"AA",x"04",x"D7",x"BE",x"AD",x"5E",x"AB",x"D0",x"0D",x"87",x"AE",x"08",x"4C",x"99",x"C1",x"AF",x"B7",x"A7",x"4A",x"EE",x"A8",x"94",x"A0",x"A9",x"27",x"5F",x"2B",x"CC",x"50",x"04",x"47",x"87",x"00",x"EF",x"D7",x"85",x"19",x"46",x"04",x"61",x"28",x"D8",x"C4",x"B9",x"FF",x"B3",x"F8",x"98",x"AD",x"5D",x"08",x"E0",x"B8",x"DE",x"DB",x"32",x"6C",x"CA",x"93",x"34",x"01",x"10",x"EA",x"00",x"90",x"B4",x"55",x"02",x"1D",x"20",x"45",x"40",x"D0",x"03",x"9D",x"DD",x"B0",x"CD",x"C8",x"41",x"26",x"1B",x"3D",x"5B",x"36",x"08",x"7D",x"5C",x"04",x"40",x"BD",x"AD",x"61",x"90",x"D1",x"07",x"5F",x"7B",x"B0",x"03",x"38",x"E9",x"20",x"60",x"48",x"FF",x"A6",x"42",x"B3",x"37",x"0D",x"56",x"FF",x"F0",x"51",x"29",x"0F",x"6F",x"7D",x"C9",x"96",x"62",x"AA",x"CA",x"DA",x"67",x"FC",x"C1",x"39",x"FB",x"29",x"8B",x"10",x"6A",x"0F",x"50",x"AD",x"09",x"B5",x"60",x"8E",x"05",x"C9",x"70",x"F0",x"01",x"3E",x"20",x"C8",x"B1",x"FB",x"48",x"BF",x"42",x"F4",x"69",x"04",x"AA",x"F5",x"97",x"2A",x"86",x"BD",x"B0",x"36",x"BA",x"64",x"18",x"C5",x"02",x"EA",x"04",x"62",x"8D",x"69",x"00",x"85",x"A6",x"5E",x"A8",x"E8",x"68",x"91",x"A5",x"E8",x"01",x"DE",x"FB",x"FA",x"FE",x"09",x"11",x"AB",x"47",x"97",x"40",x"53",x"2F",x"AC",x"C6",x"41",x"6A",x"4E",x"A8",x"30",x"D0",x"B9",x"82",x"4E",x"80",x"D6",x"D8",x"67",x"7F",x"2A",x"EC",x"0D",x"B2",x"EE",x"26",x"67",x"08",x"85",x"0E",x"DD",x"49",x"58",x"73",x"EA",x"2F",x"75",x"ED",x"09",x"5B",x"09",x"03",x"6D",x"8D",x"18",x"D4",x"CA",x"8E",x"7E",x"45",x"07",x"B3",x"4D",x"11",x"3F",x"75",x"02",x"DD",x"5D",x"E5",x"01",x"EB",x"2F",x"85",x"00",x"E8",x"25",x"B5",x"04",x"40",x"DE",x"05",x"2A",x"A9",x"81",x"5D",x"0D",x"CF",x"C8",x"FD",x"FC",x"92",x"11",x"F5",x"FA",x"E8",x"F9",x"84",x"09",x"B0",x"F5",x"C1",x"6C",x"60",x"2F",x"2C",x"3F",x"01",x"C7",x"E0",x"FF",x"0C",x"92",x"BC",x"1B",x"DE",x"0E",x"52",x"D6",x"16",x"01",x"46",x"28",x"AA",x"D6",x"5A",x"AF",x"E1",x"32",x"2A",x"F1",x"BC",x"10",x"32",x"2A",x"A3",x"31",x"D8",x"85",x"A2",x"50",x"11",x"92",x"A1",x"2A",x"1F",x"10",x"C2",x"04",x"11",x"21",x"20",x"00",x"40",x"0A",x"CA",x"BB",x"55",x"D1",x"F4",x"AE",x"9B",x"DD",x"D7",x"6A",x"0B",x"AA",x"2F",x"33",x"13",x"F3",x"EC",x"E0",x"F9",x"5F",x"47",x"39",x"D7",x"6A",x"4F",x"D9",x"4B",x"A0",x"62",x"62",x"59",x"85",x"79",x"C7",x"81",x"9F",x"78",x"B5",x"B8",x"CA",x"FE",x"FA",x"8B",x"A2",x"BB",x"2B",x"2A",x"DD",x"40",x"03",x"E8",x"E0",x"B0",x"7E",x"F5",x"ED",x"A5",x"27",x"44",x"D6",x"0D",x"A6",x"F8",x"07",x"AD",x"2E",x"76",x"61",x"15",x"D0",x"A2",x"0F",x"BE",x"D3",x"EA",x"E4",x"90",x"A0",x"DE",x"B0",x"7B",x"C0",x"D0",x"EF",x"E0",x"15",x"D1",x"DD",x"E3",x"AA",x"93",x"90",x"7B",x"A0",x"B0",x"EF",x"C0",x"D0",x"BD",x"E0",x"57",x"04",x"D2",x"B7",x"BD",x"F3",x"32",x"80",x"AF",x"90",x"F7",x"A0",x"B0",x"DE",x"C0",x"3B",x"E6",x"E0",x"BA",x"42",x"9D",x"55",x"D3",x"CA",x"10",x"AC",x"9F",x"12",x"3B",x"49",x"C8",x"BB",x"89",x"09",x"F0",x"5D",x"4B",x"25",x"B4",x"6B",x"D0",x"5C",x"B5",x"FE",x"AB",x"54",x"33",x"59",x"40",x"FF",x"D7",x"99",x"A7",x"A9",x"18",x"E6",x"72",x"D0",x"D4",x"87",x"68",x"70",x"84",x"AD",x"1B",x"D6",x"EE",x"DD",x"27",x"61",x"16",x"60",x"D8",x"DE",x"08",x"48",x"DA",x"5A",x"DB",x"A5",x"47",x"D3",x"FF",x"87",x"43",x"93",x"93",x"AC",x"49",x"3C",x"CD",x"93",x"D0",x"37",x"2D",x"5E",x"AA",x"15",x"72",x"71",x"1C",x"50",x"0A",x"AA",x"81",x"AE",x"62",x"BD",x"AA",x"82",x"57",x"85",x"AF",x"A0",x"1D",x"B1",x"AE",x"20",x"D2",x"FF",x"30",x"97",x"99",x"C0",x"07",x"EE",x"88",x"10",x"F3",x"EE",x"2F",x"CC",x"65",x"C9",x"03",x"36",x"23",x"63",x"87",x"09",x"38",x"ED",x"29",x"A9",x"8C",x"CE",x"28",x"5E",x"13",x"E9",x"AF",x"D6",x"29",x"AD",x"CE",x"50",x"D4",x"2D",x"10",x"AD",x"26",x"F5",x"5E",x"55",x"BB",x"6A",x"08",x"20",x"1C",x"15",x"3D",x"89",x"57",x"0D",x"A5",x"A7",x"F0",x"F9",x"17",x"AD",x"0B",x"49",x"EB",x"ED",x"CC",x"28",x"B1",x"CB",x"29",x"7F",x"AE",x"27",x"FA",x"A4",x"09",x"80",x"91",x"A8",x"A0",x"00",x"FC",x"22",x"99",x"0C",x"AD",x"5B",x"AD",x"02",x"AE",x"49",x"FF",x"8D",x"1D",x"DE",x"06",x"CE",x"DA",x"03",x"45",x"8C",x"01",x"DC",x"20",x"EE",x"35",x"7F",x"19",x"5D",x"57",x"30",x"1D",x"04",x"47",x"EF",x"3A",x"18",x"42",x"C9",x"6F",x"A8",x"8A",x"6D",x"0A",x"6F",x"2F",x"ED",x"B7",x"6C",x"15",x"16",x"5E",x"AE",x"A9",x"34",x"9B",x"EB",x"ED",x"6E",x"D9",x"19",x"1A",x"BC",x"09",x"F7",x"0A",x"16",x"1D",x"DA",x"3B",x"AD",x"1A",x"D4",x"38",x"2A",x"52",x"67",x"02",x"29",x"7E",x"AC",x"F7",x"63",x"20",x"C6",x"35",x"8C",x"05",x"9F",x"90",x"52",x"0A",x"48",x"F5",x"8A",x"2A",x"AA",x"68",x"8D",x"9F",x"8C",x"C7",x"71",x"A8",x"8E",x"F6",x"84",x"E3",x"78",x"79",x"AA",x"CC",x"ED",x"DF",x"32",x"09",x"A5",x"17",x"F5",x"18",x"B2",x"C9",x"10",x"35",x"8A",x"EE",x"CC",x"ED",x"6F",x"30",x"06",x"D9",x"AC",x"1B",x"4F",x"AE",x"1C",x"8C",x"57",x"60",x"8E",x"6D",x"B1",x"1B",x"31",x"35",x"98",x"20",x"4D",x"36",x"FD",x"2C",x"14",x"6D",x"AE",x"24",x"25",x"BA",x"16",x"BD",x"DC",x"FB",x"D6",x"7A",x"FA",x"68",x"28",x"40",x"7F",x"49",x"0D",x"4D",x"CB",x"CD",x"A4",x"96",x"96",x"57",x"5A",x"ED",x"8E",x"AE",x"B4",x"F0",x"0D",x"C8",x"09",x"86",x"0E",x"98",x"46",x"40",x"DB",x"0A",x"12",x"BC",x"09",x"F7",x"11",x"7B",x"DE",x"34",x"07",x"A3",x"56",x"CA",x"AC",x"D0",x"08",x"3D",x"CD",x"A9",x"F0",x"3A",x"9D",x"A4",x"72",x"ED",x"47",x"C9",x"48",x"F2",x"10",x"0F",x"27",x"18",x"10",x"E2",x"68",x"29",x"80",x"74",x"D6",x"4D",x"A5",x"D0",x"0F",x"ED",x"0C",x"3A",x"86",x"EF",x"0B",x"AA",x"99",x"BA",x"4C",x"C5",x"35",x"7B",x"06",x"08",x"BD",x"4C",x"8C",x"AD",x"8D",x"B1",x"C8",x"ED",x"21",x"58",x"EB",x"3F",x"B0",x"3E",x"00",x"42",x"C9",x"C0",x"90",x"07",x"7B",x"43",x"A2",x"FF",x"38",x"3E",x"AC",x"22",x"3D",x"8A",x"18",x"60",x"FD",x"48",x"CD",x"9A",x"31",x"20",x"25",x"2B",x"10",x"5C",x"1F",x"8C",x"86",x"D0",x"0C",x"DC",x"A2",x"29",x"EC",x"F0",x"05",x"A9",x"E8",x"82",x"20",x"F6",x"1D",x"D6",x"1E",x"AC",x"34",x"11",x"18",x"6F",x"12",x"F1",x"C9",x"60",x"5A",x"A1",x"F8",x"C9",x"00",x"F0",x"F6",x"11",x"09",x"91",x"01",x"09",x"B1",x"12",x"29",x"FE",x"BB",x"10",x"D6",x"18",x"6C",x"13",x"2D",x"9B",x"C6",x"2A",x"14",x"56",x"69",x"94",x"35",x"24",x"2A",x"AD",x"23",x"32",x"8D",x"01",x"FA",x"D0",x"60",x"47",x"15",x"A0",x"04",x"F0",x"05",x"58",x"06",x"08",x"10",x"07",x"00",x"28",x"50",x"78",x"A0",x"C8",x"F0",x"FF",x"18",x"40",x"68",x"90",x"B8",x"E0",x"08",x"30",x"FF",x"58",x"80",x"A8",x"D0",x"F8",x"20",x"48",x"70",x"FF",x"98",x"C0",x"17",x"D8",x"1E",x"D9",x"0B",x"DA",x"01",x"DB",x"22",x"91",x"D0",x"84",x"33",x"2B",x"22",x"1A",x"91",x"88",x"D0",x"5E",x"85",x"BB",x"B3",x"22",x"22",x"12",x"19",x"10",x"08",x"02",x"21",x"91",x"91",x"08",x"B9",x"5E",x"22",x"99",x"E6",x"07",x"88",x"D0",x"F7",x"18",x"AA",x"98",x"29",x"0F",x"99",x"68",x"03",x"F0",x"0C",x"8A",x"79",x"67",x"03",x"99",x"68",x"03",x"A5",x"9F",x"79",x"9B",x"03",x"99",x"9C",x"03",x"A9",x"01",x"85",x"9F",x"A9",x"78",x"20",x"00",x"01",x"4A",x"AA",x"F0",x"09",x"08",x"06",x"9F",x"38",x"6A",x"CA",x"D0",x"F9",x"28",x"6A",x"99",x"34",x"03",x"30",x"05",x"A5",x"9F",x"86",x"9F",x"24",x"8A",x"C8",x"C0",x"34",x"D0",x"C1",x"A0",x"C8",x"8A",x"4C",x"9C",x"01",x"22",x"00",x"36",x"69",x"80",x"0A",x"10",x"0F",x"06",x"FD",x"D0",x"08",x"48",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"68",x"2A",x"30",x"F1",x"70",x"01",x"60",x"38",x"85",x"A7",x"AD",x"29",x"01",x"D0",x"06",x"CE",x"2A",x"01",x"8E",x"E7",x"DB",x"CE",x"29",x"01",x"AD",x"68",x"21",x"60",x"20",x"1A",x"01",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"66",x"A8",x"CA",x"06",x"FD",x"D0",x"06",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"E8",x"90",x"F3",x"F0",x"E1",x"E0",x"11",x"B0",x"51",x"BD",x"33",x"03",x"20",x"00",x"01",x"7D",x"67",x"03",x"85",x"9E",x"AA",x"24",x"A8",x"10",x"09",x"70",x"07",x"A9",x"00",x"20",x"05",x"01",x"D0",x"25",x"A9",x"F1",x"E0",x"03",x"B0",x"03",x"BD",x"A2",x"01",x"B8",x"20",x"05",x"01",x"18",x"AA",x"BD",x"34",x"03",x"20",x"00",x"01",x"7D",x"68",x"03",x"85",x"AE",x"A5",x"A7",x"7D",x"9C",x"03",x"65",x"FF",x"85",x"AF",x"A6",x"9E",x"B1",x"AE",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"CA",x"D0",x"F1",x"86",x"A7",x"F0",x"99",x"4C",x"0D",x"08",x"CC",x"F2",x"01",x"00",x"0B",x"08",x"0A",x"7C",x"9E",x"32",x"30",x"FA",x"31",x"D3",x"A5",x"4C",x"22",x"11",x"5C",x"52",x"E8",x"50",x"53",x"09",x"45",x"9B",x"2E",x"53",x"41",x"A4",x"D2",x"3D",x"43",x"4F",x"4E",x"46",x"49",x"7E",x"55",x"52",x"D4",x"20",x"A2",x"4D",x"45",x"47",x"41",x"5F",x"B9",x"BA",x"51",x"0C",x"36",x"F5",x"13",x"50",x"52",x"4F",x"50",x"2E",x"4D",x"36",x"35",x"55",x"2E",x"4E",x"41",x"4D",x"45",x"3D",x"43",x"4F",x"4E",x"46",x"49",x"47",x"55",x"52",x"45",x"20",x"4D",x"45",x"47",x"41",x"36",x"35",x"4D",x"36",x"35",x"55",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"46",x"44",x"49",x"53",x"4B",x"2B",x"46",x"4F",x"52",x"4D",x"41",x"54",x"20",x"55",x"54",x"49",x"4C",x"49",x"54",x"59",x"00",x"00",x"00",x"00",x"00",x"E8",x"32",x"0D",x"08",x"30",x"23",x"44",x"56",x"01",x"08",x"0B",x"08",x"37",x"01",x"9E",x"32",x"30",x"36",x"31",x"00",x"00",x"00",x"BA",x"BD",x"DF",x"39",x"9D",x"FC",x"00",x"CA",x"D0",x"F7",x"A0",x"35",x"4C",x"91",x"39",x"90",x"76",x"D7",x"9A",x"AE",x"75",x"E9",x"79",x"86",x"3F",x"60",x"05",x"A2",x"A1",x"E8",x"E9",x"01",x"FA",x"08",x"23",x"D8",x"B7",x"37",x"47",x"08",x"1F",x"3D",x"32",x"CB",x"5F",x"E8",x"7C",x"F1",x"4D",x"83",x"B3",x"49",x"7D",x"DE",x"4A",x"7A",x"CB",x"4B",x"AB",x"A6",x"B0",x"4C",x"B5",x"9C",x"63",x"E6",x"A1",x"8D",x"67",x"F8",x"50",x"8E",x"68",x"9C",x"30",x"69",x"EE",x"0F",x"9D",x"51",x"6A",x"3C",x"14",x"8D",x"6B",x"1F",x"8E",x"8A",x"6C",x"13",x"C6",x"6D",x"0B",x"BD",x"38",x"6E",x"8A",x"84",x"0C",x"B6",x"53",x"1E",x"8D",x"8A",x"57",x"0F",x"8E",x"58",x"C5",x"09",x"A3",x"65",x"59",x"5F",x"20",x"9C",x"15",x"5A",x"B3",x"30",x"8D",x"5B",x"17",x"8E",x"5C",x"E6",x"04",x"C4",x"5D",x"DA",x"78",x"AA",x"87",x"2B",x"5E",x"95",x"6A",x"10",x"18",x"42",x"A3",x"93",x"C4",x"61",x"59",x"77",x"17",x"91",x"02",x"D2",x"01",x"8A",x"14",x"02",x"8B",x"9E",x"09",x"20",x"F0",x"0B",x"C1",x"5A",x"05",x"90",x"42",x"FF",x"C3",x"CA",x"B2",x"E8",x"70",x"40",x"E6",x"34",x"11",x"24",x"9C",x"EA",x"EB",x"81",x"8E",x"71",x"05",x"3E",x"C8",x"B2",x"20",x"70",x"89",x"05",x"E5",x"1A",x"8B",x"F2",x"8B",x"52",x"B2",x"61",x"F2",x"11",x"1F",x"4D",x"72",x"75",x"AB",x"54",x"76",x"41",x"6F",x"77",x"15",x"61",x"8D",x"78",x"7B",x"09",x"FB",x"9B",x"38",x"84",x"11",x"BC",x"90",x"2F",x"F2",x"24",x"06",x"C8",x"48",x"03",x"2F",x"73",x"DC",x"B2",x"C8",x"02",x"0A",x"58",x"81",x"66",x"6A",x"3D",x"12",x"DB",x"B6",x"C2",x"59",x"03",x"7D",x"EB",x"55",x"8F",x"AD",x"A9",x"AA",x"D4",x"8D",x"90",x"7B",x"11",x"4F",x"7E",x"22",x"0C",x"E0",x"32",x"E3",x"2D",x"83",x"63",x"DA",x"9E",x"05",x"BC",x"AB",x"68",x"D6",x"4B",x"36",x"FB",x"1E",x"F1",x"3C",x"0B",x"D8",x"EA",x"BA",x"50",x"79",x"BC",x"8C",x"0A",x"08",x"05",x"E2",x"41",x"68",x"21",x"C8",x"76",x"36",x"0B",x"03",x"BA",x"23",x"92",x"1F",x"0F",x"8F",x"E2",x"EB",x"3A",x"8E",x"39",x"69",x"46",x"F8",x"20",x"47",x"F8",x"07",x"6F",x"B9",x"53",x"EC",x"15",x"78",x"33",x"65",x"D3",x"BD",x"83",x"FA",x"80",x"82",x"B4",x"5A",x"AB",x"29",x"1A",x"00",x"D2",x"15",x"2D",x"47",x"0C",x"FB",x"01",x"E5",x"0F",x"68",x"14",x"8A",x"F6",x"A8",x"FC",x"41",x"CD",x"E0",x"81",x"F0",x"FE",x"47",x"79",x"95",x"83",x"F0",x"0D",x"A4",x"DC",x"3F",x"80",x"64",x"12",x"15",x"98",x"AC",x"5A",x"C4",x"55",x"CA",x"4E",x"C5",x"77",x"0D",x"1B",x"07",x"AC",x"B9",x"37",x"FE",x"78",x"37",x"62",x"9C",x"A4",x"C4",x"2B",x"78",x"3E",x"B7",x"B4",x"CC",x"20",x"C9",x"4A",x"FF",x"70",x"F7",x"78",x"10",x"A0",x"C2",x"1B",x"CE",x"8B",x"01",x"1A",x"F5",x"D1",x"FA",x"83",x"D4",x"EC",x"12",x"27",x"2D",x"6E",x"D1",x"A9",x"26",x"D2",x"CB",x"A1",x"D2",x"D8",x"A9",x"2F",x"94",x"AF",x"D7",x"B6",x"F3",x"32",x"51",x"CD",x"CE",x"EF",x"CF",x"59",x"34",x"C2",x"A8",x"DE",x"0D",x"FC",x"F8",x"35",x"0D",x"CE",x"67",x"FF",x"DC",x"D3",x"E4",x"D4",x"3D",x"D5",x"66",x"C7",x"D6",x"7C",x"E7",x"8B",x"5A",x"71",x"D9",x"33",x"33",x"E1",x"3E",x"70",x"05",x"90",x"A6",x"13",x"42",x"29",x"A9",x"A1",x"61",x"EF",x"0F",x"58",x"00",x"22",x"72",x"3F",x"57",x"E0",x"34",x"A6",x"91",x"9D",x"D3",x"E8",x"E7",x"04",x"79",x"56",x"C7",x"B0",x"A6",x"18",x"88",x"ED",x"AA",x"CF",x"13",x"78",x"C8",x"00",x"7F",x"8F",x"0F",x"07",x"F0",x"7B",x"05",x"BD",x"10",x"6B",x"43",x"6A",x"91",x"8D",x"EF",x"14",x"4C",x"00",x"18",x"1F",x"1C",x"3E",x"1E",x"CC",x"A6",x"A9",x"40",x"28",x"01",x"24",x"AC",x"39",x"28",x"AA",x"3F",x"35",x"EA",x"42",x"9C",x"40",x"C7",x"3D",x"28",x"E5",x"0F",x"79",x"E9",x"2C",x"5E",x"C6",x"2B",x"84",x"13",x"A3",x"A9",x"2E",x"DD",x"E9",x"60",x"48",x"EA",x"50",x"A2",x"0B",x"E2",x"04",x"CD",x"A2",x"18",x"8D",x"EB",x"08",x"D3",x"D2",x"BC",x"7C",x"C9",x"16",x"A4",x"57",x"14",x"3B",x"F1",x"40",x"08",x"4C",x"42",x"91",x"A6",x"92",x"EC",x"80",x"93",x"AD",x"0C",x"94",x"53",x"9C",x"95",x"9A",x"32",x"22",x"96",x"A9",x"A9",x"41",x"97",x"EB",x"98",x"99",x"BD",x"9A",x"F7",x"9B",x"4A",x"8D",x"9C",x"79",x"1F",x"E6",x"9E",x"A2",x"73",x"E0",x"5C",x"79",x"82",x"A1",x"53",x"79",x"D2",x"00",x"B3",x"0A",x"19",x"E6",x"01",x"8D",x"B1",x"79",x"60",x"F9",x"47",x"51",x"8B",x"26",x"F5",x"4F",x"B9",x"FB",x"73",x"F3",x"51",x"D6",x"2B",x"51",x"5D",x"1E",x"6F",x"BE",x"5C",x"51",x"82",x"DD",x"B4",x"9C",x"1B",x"2A",x"07",x"9C",x"D1",x"F1",x"05",x"E2",x"1C",x"03",x"74",x"39",x"10",x"5E",x"61",x"06",x"02",x"E1",x"06",x"04",x"7C",x"03",x"0C",x"AF",x"01",x"06",x"F5",x"04",x"B1",x"07",x"81",x"05",x"8F",x"2C",x"06",x"08",x"A7",x"4B",x"02",x"79",x"A4",x"79",x"9F",x"2C",x"33",x"0A",x"06",x"36",x"31",x"45",x"01",x"E3",x"A5",x"29",x"70",x"5A",x"2F",x"17",x"7D",x"BE",x"E3",x"0F",x"B5",x"0E",x"AB",x"5D",x"09",x"2F",x"7C",x"5A",x"89",x"AC",x"80",x"5C",x"DB",x"5C",x"21",x"47",x"2E",x"04",x"1E",x"70",x"1A",x"08",x"88",x"8A",x"01",x"B3",x"91",x"BC",x"74",x"6A",x"41",x"50",x"56",x"5F",x"E0",x"EB",x"1E",x"0C",x"1F",x"64",x"E0",x"AB",x"67",x"09",x"80",x"CB",x"6F",x"67",x"3F",x"43",x"04",x"29",x"5D",x"61",x"9A",x"05",x"7F",x"C3",x"E2",x"4F",x"11",x"2A",x"DA",x"29",x"80",x"26",x"0E",x"5E",x"A8",x"16",x"6A",x"5A",x"0C",x"83",x"0F",x"14",x"27",x"10",x"C0",x"13",x"87",x"13",x"13",x"E0",x"12",x"C3",x"0C",x"1B",x"F0",x"0D",x"A1",x"7B",x"86",x"06",x"2A",x"1F",x"0F",x"EE",x"18",x"5E",x"0B",x"2E",x"7C",x"0E",x"B8",x"4D",x"36",x"7C",x"15",x"B8",x"3E",x"C6",x"94",x"31",x"E8",x"33",x"91",x"0F",x"0D",x"7A",x"23",x"79",x"97",x"A1",x"8A",x"66",x"04",x"1E",x"89",x"4C",x"C5",x"79",x"A1",x"35",x"99",x"ED",x"1D",x"39",x"5D",x"A4",x"04",x"F3",x"EE",x"3F",x"38",x"5F",x"21",x"C8",x"5A",x"38",x"B0",x"F2",x"F2",x"14",x"8A",x"C1",x"94",x"A3",x"A0",x"66",x"D4",x"E3",x"E0",x"F2",x"62",x"E7",x"09",x"1A",x"B2",x"D0",x"7E",x"4B",x"7D",x"8F",x"A8",x"64",x"55",x"D0",x"07",x"AD",x"90",x"7B",x"C9",x"88",x"FF",x"2C",x"44",x"B5",x"71",x"3A",x"0E",x"18",x"C9",x"A9",x"7D",x"B5",x"41",x"85",x"04",x"B0",x"F3",x"3F",x"20",x"2E",x"0F",x"E5",x"3B",x"34",x"F0",x"35",x"85",x"FB",x"9F",x"62",x"AD",x"29",x"D6",x"8D",x"5B",x"BF",x"FC",x"6B",x"7C",x"0C",x"72",x"41",x"80",x"80",x"0A",x"76",x"9B",x"5C",x"68",x"99",x"A3",x"CF",x"B3",x"85",x"50",x"9C",x"CB",x"73",x"62",x"73",x"6B",x"37",x"47",x"64",x"4E",x"39",x"60",x"CA",x"E9",x"61",x"02",x"1C",x"F7",x"CC",x"07",x"39",x"80",x"1B",x"FB",x"3C",x"86",x"E9",x"BC",x"00",x"8C",x"9F",x"F1",x"00",x"8A",x"6E",x"E5",x"FD",x"49",x"30",x"0F",x"13",x"B1",x"20",x"A0",x"5F",x"60",x"67",x"60",x"1B",x"C8",x"1D",x"E9",x"91",x"64",x"2B",x"82",x"A8",x"B9",x"19",x"E7",x"0A",x"95",x"64",x"17",x"DF",x"10",x"CB",x"A7",x"02",x"9D",x"2F",x"1D",x"A0",x"A8",x"B9",x"49",x"F6",x"75",x"B0",x"97",x"E5",x"10",x"CC",x"45",x"50",x"B8",x"93",x"E4",x"B6",x"9A",x"09",x"C5",x"04",x"7E",x"E2",x"C5",x"CB",x"9A",x"B2",x"35",x"06",x"EB",x"B6",x"78",x"74",x"15",x"99",x"99",x"85",x"5C",x"6F",x"41",x"82",x"62",x"60",x"00",x"E1",x"DE",x"65",x"79",x"B9",x"63",x"11",x"B2",x"41",x"B8",x"B9",x"24",x"CF",x"02",x"1F",x"A4",x"57",x"86",x"80",x"88",x"3C",x"A1",x"3A",x"B2",x"C5",x"1C",x"99",x"03",x"E1",x"C4",x"13",x"23",x"F1",x"04",x"B2",x"CB",x"D0",x"D8",x"D5",x"AC",x"51",x"77",x"AD",x"03",x"7A",x"E0",x"13",x"A2",x"8B",x"F9",x"3D",x"82",x"FD",x"40",x"03",x"45",x"26",x"05",x"07",x"48",x"AD",x"90",x"06",x"A4",x"56",x"48",x"05",x"4A",x"AD",x"04",x"7A",x"84",x"5F",x"21",x"B3",x"90",x"E6",x"2A",x"4F",x"00",x"57",x"13",x"1B",x"EE",x"E0",x"19",x"05",x"4F",x"D7",x"13",x"F0",x"1C",x"F0",x"B7",x"06",x"D0",x"05",x"AA",x"1A",x"3C",x"0D",x"68",x"25",x"CF",x"71",x"CF",x"B8",x"E0",x"87",x"35",x"A9",x"40",x"EF",x"E3",x"2A",x"20",x"55",x"2C",x"7D",x"3D",x"41",x"32",x"AC",x"1C",x"0D",x"2F",x"80",x"F9",x"90",x"6F",x"B6",x"75",x"03",x"A0",x"24",x"20",x"63",x"65",x"16",x"1F",x"23",x"05",x"D2",x"50",x"DD",x"02",x"8D",x"BA",x"2D",x"C6",x"1B",x"C3",x"26",x"85",x"9E",x"95",x"F2",x"04",x"44",x"88",x"F9",x"2B",x"AD",x"0E",x"E0",x"4E",x"9D",x"20",x"30",x"81",x"87",x"B6",x"41",x"73",x"A3",x"30",x"70",x"04",x"39",x"1D",x"CD",x"31",x"B1",x"8A",x"21",x"53",x"75",x"01",x"64",x"EC",x"55",x"02",x"87",x"6E",x"A0",x"5F",x"B2",x"C4",x"2B",x"5F",x"8A",x"A1",x"5E",x"2C",x"85",x"42",x"5D",x"4A",x"AD",x"5C",x"77",x"B2",x"27",x"DE",x"BD",x"1C",x"6E",x"94",x"EA",x"93",x"29",x"63",x"92",x"4A",x"A9",x"5E",x"B4",x"4F",x"36",x"A9",x"37",x"F7",x"38",x"7C",x"9D",x"19",x"5F",x"98",x"15",x"43",x"97",x"B4",x"14",x"2A",x"96",x"52",x"7A",x"B5",x"79",x"3A",x"AD",x"3B",x"F7",x"3C",x"32",x"D4",x"19",x"F1",x"98",x"54",x"D9",x"AA",x"61",x"D9",x"24",x"47",x"01",x"4A",x"AB",x"6B",x"04",x"3B",x"1A",x"D2",x"B3",x"0F",x"18",x"E3",x"19",x"07",x"16",x"4B",x"16",x"80",x"F0",x"12",x"9A",x"78",x"47",x"F9",x"4B",x"20",x"09",x"E5",x"89",x"E4",x"0F",x"F8",x"CC",x"F4",x"20",x"99",x"42",x"7D",x"79",x"B4",x"73",x"A9",x"EB",x"9B",x"01",x"EB",x"4D",x"7D",x"88",x"AB",x"72",x"F7",x"22",x"C5",x"F0",x"81",x"B7",x"F4",x"4B",x"DD",x"8C",x"0E",x"82",x"50",x"4F",x"8F",x"AC",x"38",x"2F",x"91",x"6C",x"A2",x"73",x"FE",x"28",x"42",x"2B",x"2D",x"7E",x"5E",x"CA",x"24",x"CC",x"C8",x"C8",x"3A",x"7F",x"D8",x"38",x"6F",x"10",x"2A",x"51",x"4F",x"0A",x"C8",x"FC",x"4F",x"63",x"87",x"EA",x"34",x"9C",x"99",x"79",x"D9",x"A9",x"F0",x"73",x"1F",x"05",x"75",x"8A",x"59",x"77",x"CB",x"32",x"A5",x"35",x"8B",x"AB",x"C5",x"9A",x"AB",x"8A",x"0E",x"C8",x"96",x"7B",x"42",x"B3",x"0C",x"77",x"22",x"6F",x"24",x"F0",x"CF",x"20",x"BC",x"7B",x"38",x"2F",x"B9",x"80",x"F0",x"96",x"29",x"37",x"7B",x"80",x"6A",x"96",x"CB",x"19",x"0C",x"40",x"2A",x"B9",x"83",x"98",x"40",x"BB",x"C2",x"0D",x"6E",x"CD",x"7B",x"A9",x"C2",x"19",x"F6",x"7C",x"3E",x"18",x"C3",x"14",x"4C",x"E0",x"23",x"3D",x"F5",x"3C",x"3C",x"3B",x"3A",x"EF",x"6A",x"44",x"68",x"F0",x"60",x"D5",x"EF",x"BD",x"35",x"E3",x"34",x"79",x"33",x"B6",x"66",x"E8",x"07",x"A7",x"4E",x"E5",x"DC",x"8D",x"4E",x"41",x"EB",x"40",x"59",x"6B",x"40",x"AD",x"56",x"AD",x"B3",x"45",x"3E",x"78",x"3F",x"40",x"CF",x"41",x"90",x"F3",x"FB",x"F7",x"01",x"78",x"97",x"EB",x"38",x"07",x"4F",x"C5",x"CD",x"85",x"58",x"D0",x"74",x"39",x"5A",x"64",x"80",x"11",x"5F",x"28",x"73",x"D8",x"EB",x"AD",x"39",x"E0",x"38",x"75",x"C9",x"6E",x"37",x"4A",x"AD",x"36",x"4B",x"8D",x"32",x"4B",x"8E",x"33",x"8B",x"BD",x"34",x"2A",x"B5",x"8D",x"35",x"5F",x"4C",x"96",x"17",x"E2",x"4C",x"8D",x"A7",x"16",x"BF",x"9B",x"4B",x"B7",x"E5",x"22",x"B9",x"2F",x"5F",x"92",x"16",x"94",x"BC",x"50",x"C7",x"AA",x"FB",x"15",x"DC",x"F0",x"EE",x"F0",x"00",x"C1",x"7B",x"85",x"19",x"01",x"80",x"B9",x"18",x"68",x"13",x"BC",x"19",x"2C",x"AE",x"48",x"A9",x"93",x"E0",x"A3",x"50",x"3F",x"95",x"B7",x"72",x"02",x"9E",x"6D",x"E0",x"08",x"1F",x"F9",x"63",x"40",x"98",x"09",x"F4",x"2D",x"0F",x"17",x"4C",x"14",x"40",x"3E",x"EC",x"6E",x"A7",x"5D",x"C4",x"9A",x"F8",x"85",x"23",x"C4",x"AA",x"29",x"DC",x"F5",x"63",x"03",x"EC",x"75",x"C1",x"7C",x"AA",x"30",x"2F",x"08",x"91",x"8D",x"91",x"1C",x"5A",x"01",x"08",x"D6",x"06",x"30",x"62",x"0E",x"A1",x"29",x"F1",x"32",x"F0",x"E1",x"4D",x"EB",x"31",x"95",x"D9",x"A5",x"CD",x"E6",x"72",x"86",x"64",x"B9",x"94",x"1A",x"B3",x"7E",x"88",x"93",x"AB",x"5D",x"52",x"BD",x"32",x"F8",x"20",x"EF",x"48",x"F2",x"B9",x"7A",x"BA",x"BB",x"4F",x"A1",x"C1",x"4C",x"CE",x"50",x"19",x"FA",x"96",x"E3",x"1C",x"F5",x"69",x"B0",x"AE",x"83",x"9D",x"82",x"8F",x"C9",x"01",x"AD",x"3C",x"B4",x"B2",x"40",x"64",x"12",x"1D",x"0E",x"51",x"C1",x"B4",x"8C",x"A0",x"B4",x"40",x"79",x"9C",x"48",x"61",x"AB",x"08",x"B7",x"A8",x"E3",x"4F",x"F7",x"1A",x"8A",x"BD",x"DB",x"4B",x"C1",x"C2",x"BD",x"C3",x"E7",x"C4",x"79",x"BC",x"BB",x"CF",x"BA",x"F3",x"B9",x"56",x"43",x"08",x"F2",x"74",x"3F",x"E3",x"F4",x"E0",x"C9",x"CA",x"BC",x"CB",x"67",x"D1",x"08",x"E0",x"03",x"3F",x"4B",x"B0",x"06",x"4D",x"24",x"8D",x"59",x"8E",x"D6",x"34",x"1D",x"E1",x"4C",x"47",x"84",x"A9",x"90",x"80",x"79",x"C7",x"71",x"57",x"7E",x"7F",x"EF",x"80",x"59",x"33",x"C2",x"AE",x"78",x"00",x"4C",x"80",x"7A",x"1E",x"5F",x"D1",x"03",x"A1",x"94",x"48",x"0C",x"0A",x"77",x"94",x"74",x"BE",x"67",x"E2",x"82",x"6A",x"94",x"1B",x"F2",x"B4",x"B6",x"D1",x"BC",x"0F",x"A9",x"5C",x"92",x"49",x"3A",x"5D",x"0C",x"CE",x"F8",x"1D",x"A3",x"DC",x"7E",x"5E",x"64",x"20",x"9F",x"CA",x"AD",x"11",x"AB",x"28",x"BE",x"38",x"3A",x"E8",x"25",x"A3",x"C5",x"1F",x"14",x"D4",x"2B",x"9B",x"3A",x"04",x"A8",x"F2",x"F1",x"8E",x"B2",x"A9",x"AD",x"92",x"E9",x"94",x"53",x"74",x"DD",x"5B",x"16",x"D2",x"B8",x"E5",x"34",x"7D",x"1E",x"A5",x"1C",x"6F",x"A0",x"D9",x"DA",x"DE",x"DB",x"73",x"87",x"53",x"89",x"6E",x"64",x"76",x"DC",x"15",x"31",x"DB",x"DA",x"CF",x"D9",x"2B",x"40",x"E0",x"C4",x"DF",x"F3",x"DE",x"DD",x"BC",x"87",x"3E",x"68",x"A3",x"1B",x"62",x"1D",x"CB",x"C4",x"3C",x"AF",x"D4",x"6D",x"9A",x"8A",x"01",x"44",x"0E",x"12",x"CC",x"47",x"1B",x"BA",x"A8",x"8A",x"B6",x"E1",x"4E",x"C1",x"8B",x"DA",x"CD",x"01",x"22",x"13",x"E0",x"A2",x"08",x"BB",x"2A",x"8E",x"D9",x"CF",x"A4",x"62",x"9C",x"64",x"12",x"EF",x"7D",x"00",x"47",x"83",x"5A",x"BD",x"A6",x"8E",x"BE",x"B4",x"D8",x"CB",x"BF",x"52",x"2F",x"47",x"E2",x"47",x"45",x"84",x"E7",x"8B",x"83",x"29",x"B7",x"29",x"8D",x"19",x"8F",x"DD",x"90",x"B3",x"68",x"84",x"CF",x"D9",x"07",x"15",x"92",x"F0",x"93",x"94",x"9E",x"45",x"23",x"C2",x"CC",x"3E",x"6B",x"A8",x"0F",x"79",x"64",x"5C",x"86",x"87",x"EF",x"88",x"A9",x"63",x"89",x"4A",x"E2",x"3C",x"EF",x"28",x"DE",x"50",x"96",x"97",x"EF",x"98",x"A9",x"B9",x"99",x"78",x"1E",x"F3",x"1E",x"E4",x"73",x"9C",x"03",x"1E",x"E0",x"72",x"1E",x"C0",x"6E",x"10",x"BA",x"AC",x"B3",x"07",x"C4",x"2C",x"04",x"B0",x"C1",x"03",x"FA",x"80",x"09",x"1C",x"20",x"31",x"17",x"0F",x"B0",x"07",x"C4",x"24",x"2E",x"EA",x"33",x"0B",x"13",x"03",x"F0",x"C7",x"EF",x"C8",x"07",x"15",x"DE",x"04",x"16",x"6C",x"8A",x"8B",x"BC",x"35",x"E3",x"41",x"09",x"29",x"0B",x"88",x"19",x"82",x"AE",x"A5",x"83",x"78",x"4D",x"B3",x"06",x"9B",x"3B",x"E1",x"57",x"A2",x"07",x"A6",x"D7",x"17",x"38",x"DE",x"ED",x"7A",x"06",x"7E",x"B4",x"17",x"4C",x"8E",x"D6",x"27",x"6D",x"05",x"6C",x"E8",x"78",x"03",x"1B",x"04",x"1B",x"64",x"2E",x"03",x"34",x"BA",x"91",x"76",x"A3",x"0A",x"00",x"A2",x"5E",x"E7",x"11",x"05",x"23",x"29",x"7B",x"82",x"6A",x"70",x"B5",x"66",x"18",x"69",x"52",x"DC",x"7C",x"02",x"B5",x"EC",x"C3",x"91",x"5E",x"38",x"1B",x"18",x"0F",x"57",x"D6",x"55",x"4A",x"14",x"A1",x"9F",x"5B",x"FF",x"D0",x"E9",x"23",x"25",x"65",x"3D",x"F8",x"D4",x"87",x"6E",x"F8",x"73",x"4D",x"AC",x"18",x"89",x"E8",x"44",x"53",x"4E",x"06",x"D3",x"D6",x"B1",x"C3",x"AE",x"CA",x"36",x"10",x"F1",x"14",x"A3",x"B2",x"6A",x"CC",x"6A",x"40",x"08",x"AE",x"6A",x"71",x"4D",x"02",x"C8",x"4D",x"26",x"A6",x"A0",x"D2",x"01",x"50",x"07",x"BA",x"15",x"35",x"B7",x"9B",x"92",x"E5",x"45",x"2F",x"66",x"50",x"FD",x"4A",x"21",x"3E",x"04",x"97",x"A2",x"F5",x"88",x"9E",x"17",x"55",x"E5",x"AF",x"5C",x"4C",x"0E",x"33",x"27",x"19",x"7D",x"EB",x"E5",x"A9",x"09",x"12",x"DC",x"2A",x"E7",x"70",x"A0",x"10",x"49",x"01",x"8F",x"3D",x"20",x"5D",x"FE",x"A8",x"09",x"3E",x"69",x"0E",x"19",x"62",x"F0",x"DE",x"0A",x"73",x"6D",x"60",x"77",x"F9",x"95",x"56",x"99",x"7D",x"70",x"85",x"2F",x"A0",x"C0",x"00",x"80",x"04",x"AA",x"EF",x"0F",x"C8",x"B9",x"BF",x"73",x"FA",x"D9",x"E1",x"7C",x"F0",x"F4",x"7F",x"01",x"B0",x"02",x"FA",x"FF",x"0B",x"53",x"F6",x"F0",x"13",x"B9",x"D2",x"18",x"62",x"08",x"86",x"EC",x"B4",x"05",x"54",x"82",x"80",x"06",x"AE",x"4C",x"BD",x"4C",x"FE",x"22",x"EE",x"7C",x"11",x"4E",x"6C",x"56",x"0C",x"A8",x"24",x"6B",x"BB",x"ED",x"A0",x"08",x"92",x"CC",x"2C",x"C4",x"03",x"F2",x"24",x"42",x"0F",x"7B",x"6A",x"5E",x"27",x"83",x"81",x"08",x"E3",x"DF",x"0D",x"22",x"61",x"D5",x"12",x"5D",x"1D",x"6B",x"95",x"C4",x"E1",x"C3",x"79",x"C2",x"C1",x"5E",x"D1",x"46",x"0C",x"9B",x"3B",x"90",x"CE",x"FA",x"5C",x"3A",x"00",x"FB",x"0E",x"F6",x"56",x"E2",x"4D",x"2E",x"03",x"4F",x"0F",x"9E",x"FD",x"34",x"E2",x"3B",x"39",x"50",x"D9",x"0E",x"79",x"E6",x"C0",x"91",x"47",x"60",x"D5",x"CF",x"70",x"62",x"34",x"F0",x"C5",x"A7",x"C0",x"8C",x"BF",x"E7",x"BE",x"79",x"BD",x"71",x"A2",x"1E",x"CC",x"F2",x"A5",x"49",x"E8",x"CE",x"6D",x"9A",x"ED",x"10",x"71",x"D0",x"E0",x"CF",x"79",x"CE",x"CD",x"DE",x"D1",x"C4",x"D2",x"6B",x"74",x"10",x"71",x"D6",x"E0",x"D5",x"79",x"D4",x"D3",x"DE",x"1F",x"D7",x"44",x"AE",x"D8",x"7C",x"E9",x"BA",x"EB",x"45",x"10",x"97",x"05",x"CC",x"D2",x"CB",x"F3",x"CA",x"C9",x"BC",x"5A",x"44",x"8D",x"3C",x"8C",x"8B",x"CF",x"8A",x"9B",x"3E",x"B8",x"09",x"45",x"0E",x"1E",x"06",x"D8",x"54",x"58",x"6E",x"13",x"81",x"80",x"9E",x"7F",x"A7",x"E3",x"7E",x"78",x"D6",x"D4",x"0A",x"56",x"12",x"01",x"FB",x"31",x"A0",x"90",x"C2",x"19",x"06",x"DC",x"92",x"28",x"B8",x"30",x"01",x"12",x"8B",x"8C",x"64",x"46",x"8E",x"63",x"11",x"35",x"01",x"F9",x"04",x"40",x"35",x"C8",x"17",x"BC",x"1C",x"A4",x"EC",x"31",x"86",x"79",x"9A",x"C9",x"7D",x"27",x"37",x"62",x"A3",x"9B",x"20",x"9F",x"CB",x"0A",x"83",x"58",x"00",x"38",x"42",x"C7",x"02",x"58",x"32",x"AF",x"08",x"B1",x"9B",x"A2",x"E1",x"B2",x"F4",x"0A",x"4D",x"C9",x"02",x"64",x"60",x"C0",x"97",x"45",x"5A",x"FF",x"70",x"0B",x"A0",x"4B",x"B0",x"10",x"A0",x"92",x"0E",x"B0",x"1C",x"54",x"2D",x"A0",x"06",x"12",x"64",x"D7",x"D1",x"73",x"00",x"BB",x"1A",x"1D",x"A0",x"7E",x"B0",x"EB",x"D0",x"63",x"00",x"BB",x"18",x"29",x"A0",x"7E",x"B0",x"EB",x"01",x"58",x"76",x"F4",x"34",x"00",x"C8",x"55",x"4C",x"64",x"C7",x"29",x"11",x"C6",x"52",x"AA",x"C5",x"7C",x"56",x"91",x"89",x"7A",x"88",x"C1",x"DE",x"87",x"A6",x"54",x"86",x"79",x"EF",x"C3",x"A6",x"AD",x"5C",x"57",x"73",x"78",x"01",x"D3",x"C1",x"EF",x"4E",x"E7",x"B4",x"5A",x"73",x"F5",x"49",x"90",x"71",x"EA",x"35",x"09",x"2C",x"13",x"08",x"1B",x"D7",x"CC",x"92",x"F8",x"72",x"66",x"34",x"90",x"55",x"79",x"2B",x"9B",x"A5",x"F0",x"22",x"A9",x"91",x"9D",x"2E",x"C7",x"73",x"0C",x"33",x"08",x"71",x"97",x"2B",x"A0",x"FF",x"C8",x"B9",x"12",x"73",x"99",x"FF",x"E1",x"7C",x"D0",x"F7",x"8F",x"43",x"8D",x"E2",x"E3",x"30",x"57",x"B9",x"90",x"EE",x"5E",x"93",x"7C",x"1A",x"5E",x"36",x"BF",x"57",x"0B",x"1C",x"28",x"B6",x"1F",x"F4",x"A1",x"44",x"F7",x"37",x"9B",x"E1",x"A2",x"7C",x"F5",x"03",x"93",x"45",x"A8",x"81",x"2D",x"AA",x"98",x"F2",x"07",x"A9",x"4A",x"71",x"C2",x"A9",x"8D",x"25",x"20",x"DA",x"BF",x"07",x"DE",x"7B",x"DE",x"11",x"20",x"93",x"15",x"A6",x"16",x"B6",x"01",x"96",x"45",x"08",x"16",x"5A",x"0A",x"12",x"43",x"92",x"A9",x"15",x"4C",x"8B",x"2A",x"91",x"CF",x"D0",x"14",x"72",x"7E",x"6F",x"AD",x"23",x"04",x"4C",x"14",x"2C",x"E9",x"AF",x"6C",x"35",x"07",x"21",x"76",x"20",x"76",x"52",x"F2",x"B0",x"BD",x"58",x"47",x"99",x"EF",x"2B",x"82",x"91",x"3A",x"35",x"E2",x"C8",x"A8",x"8E",x"0A",x"88",x"DC",x"10",x"FC",x"6A",x"32",x"FF",x"48",x"68",x"BA",x"1E",x"AA",x"8D",x"BF",x"0B",x"B3",x"64",x"0B",x"E7",x"D1",x"30",x"55",x"CE",x"2C",x"E4",x"0B",x"D0",x"08",x"C5",x"0A",x"F0",x"09",x"FF",x"0B",x"2C",x"2C",x"0C",x"E3",x"44",x"08",x"D9",x"B0",x"8E",x"B4",x"78",x"73",x"F0",x"0D",x"E2",x"29",x"07",x"4B",x"7C",x"15",x"A7",x"57",x"5F",x"87",x"37",x"6D",x"AF",x"0C",x"CA",x"14",x"55",x"AA",x"64",x"79",x"57",x"5C",x"76",x"D2",x"2D",x"9A",x"61",x"3B",x"00",x"17",x"29",x"66",x"72",x"B5",x"51",x"5A",x"50",x"31",x"6F",x"A2",x"6D",x"80",x"0F",x"BF",x"59",x"AE",x"76",x"AE",x"6F",x"35",x"AB",x"F3",x"42",x"73",x"D5",x"93",x"A9",x"37",x"20",x"E3",x"C4",x"34",x"97",x"77",x"BA",x"D0",x"02",x"80",x"FE",x"5F",x"31",x"70",x"EB",x"01",x"96",x"39",x"FC",x"3F",x"30",x"3F",x"B2",x"E9",x"3E",x"5B",x"4C",x"0A",x"1A",x"5E",x"47",x"09",x"53",x"8D",x"2F",x"D0",x"F3",x"69",x"CA",x"17",x"7B",x"63",x"56",x"58",x"1B",x"08",x"19",x"20",x"35",x"1B",x"69",x"87",x"D0",x"7C",x"78",x"20",x"78",x"F0",x"70",x"59",x"8A",x"5B",x"A7",x"2D",x"5A",x"53",x"35",x"6B",x"50",x"04",x"B9",x"D8",x"68",x"8D",x"2E",x"54",x"A9",x"04",x"C0",x"E3",x"18",x"10",x"1D",x"60",x"29",x"DC",x"28",x"F8",x"92",x"33",x"56",x"C5",x"A4",x"58",x"5A",x"67",x"60",x"A1",x"23",x"9C",x"04",x"CB",x"04",x"1A",x"A0",x"54",x"59",x"B0",x"A1",x"E3",x"D4",x"83",x"C3",x"43",x"E2",x"58",x"0E",x"CC",x"76",x"A9",x"81",x"8B",x"70",x"58",x"22",x"64",x"40",x"54",x"3D",x"E1",x"01",x"83",x"33",x"5A",x"57",x"82",x"8C",x"58",x"76",x"31",x"AC",x"0C",x"B6",x"8D",x"D6",x"09",x"40",x"56",x"10",x"59",x"70",x"64",x"16",x"05",x"B8",x"0F",x"78",x"05",x"36",x"05",x"10",x"BC",x"06",x"0A",x"E8",x"54",x"70",x"0B",x"C6",x"4E",x"4A",x"6D",x"BA",x"4F",x"EA",x"50",x"B2",x"1A",x"A3",x"51",x"F5",x"68",x"B6",x"B4",x"40",x"52",x"2D",x"53",x"96",x"A9",x"03",x"FA",x"54",x"A9",x"9C",x"5D",x"34",x"2B",x"56",x"9E",x"71",x"55",x"CD",x"C8",x"9C",x"58",x"E9",x"90",x"D4",x"57",x"92",x"23",x"F7",x"83",x"BC",x"8A",x"20",x"E8",x"64",x"F1",x"8D",x"5A",x"3F",x"5B",x"DA",x"45",x"01",x"29",x"7F",x"DA",x"8D",x"D9",x"96",x"D0",x"70",x"E4",x"90",x"19",x"B8",x"06",x"3E",x"A6",x"33",x"E0",x"58",x"66",x"E5",x"82",x"BA",x"0C",x"5C",x"2C",x"DD",x"09",x"2F",x"5D",x"69",x"51",x"8C",x"02",x"2A",x"9C",x"04",x"4D",x"66",x"F9",x"8E",x"01",x"4D",x"A9",x"4E",x"8D",x"05",x"D7",x"7D",x"FE",x"F2",x"75",x"CC",x"E5",x"A7",x"E0",x"92",x"31",x"8E",x"ED",x"18",x"B3",x"D0",x"AD",x"73",x"56",x"29",x"FC",x"76",x"01",x"B9",x"20",x"00",x"45",x"AD",x"31",x"1B",x"09",x"03",x"76",x"DA",x"5A",x"02",x"DD",x"9C",x"20",x"7F",x"06",x"21",x"2B",x"D5",x"C9",x"8D",x"16",x"D0",x"7A",x"18",x"03",x"85",x"18",x"F9",x"68",x"19",x"16",x"4C",x"21",x"B1",x"73",x"5B",x"D2",x"8C",x"24",x"2D",x"13",x"0F",x"51",x"36",x"07",x"CA",x"D0",x"2A",x"44",x"41",x"66",x"08",x"4A",x"AE",x"09",x"56",x"1F",x"A0",x"3C",x"53",x"00",x"CA",x"C4",x"0A",x"88",x"91",x"4D",x"08",x"25",x"7B",x"26",x"7A",x"78",x"4A",x"B1",x"8E",x"A5",x"B2",x"B3",x"EF",x"B4",x"95",x"9C",x"B5",x"78",x"7E",x"7E",x"0B",x"B6",x"1A",x"02",x"7C",x"5A",x"F7",x"F6",x"B6",x"A7",x"54",x"35",x"4B",x"54",x"C4",x"54",x"48",x"03",x"17",x"D4",x"A4",x"8E",x"9C",x"1D",x"E0",x"5B",x"70",x"A9",x"F1",x"D4",x"6F",x"92",x"F1",x"D4",x"6E",x"92",x"AD",x"6D",x"D2",x"DC",x"D3",x"12",x"92",x"97",x"45",x"48",x"5B",x"51",x"AA",x"A8",x"5A",x"80",x"88",x"42",x"EC",x"50",x"20",x"E2",x"5B",x"68",x"28",x"33",x"B9",x"38",x"0F",x"EE",x"63",x"60",x"06",x"13",x"C6",x"0D",x"B1",x"65",x"27",x"72",x"C3",x"01",x"BB",x"10",x"26",x"96",x"BD",x"89",x"EA",x"B3",x"05",x"B1",x"88",x"1D",x"47",x"8E",x"51",x"A2",x"C1",x"A5",x"9A",x"8A",x"CA",x"24",x"D4",x"7E",x"B0",x"E8",x"80",x"56",x"C4",x"AB",x"E7",x"01",x"40",x"79",x"07",x"A6",x"99",x"10",x"92",x"9C",x"D9",x"A2",x"53",x"02",x"EB",x"EE",x"40",x"F2",x"0A",x"04",x"2E",x"04",x"10",x"E8",x"79",x"80",x"7C",x"50",x"D1",x"3E",x"AA",x"88",x"84",x"DD",x"DA",x"A8",x"03",x"2D",x"99",x"23",x"A3",x"FD",x"58",x"06",x"20",x"8C",x"71",x"A4",x"00",x"59",x"07",x"90",x"77",x"D1",x"81",x"64",x"2A",x"95",x"6E",x"D2",x"81",x"62",x"58",x"E5",x"91",x"78",x"3F",x"84",x"C2",x"0C",x"B0",x"9E",x"39",x"23",x"93",x"2F",x"92",x"20",x"FB",x"60",x"4E",x"A8",x"3C",x"E7",x"C4",x"C4",x"18",x"75",x"0D",x"AC",x"97",x"8D",x"5C",x"32",x"E1",x"36",x"EC",x"9C",x"4B",x"67",x"B7",x"10",x"B4",x"B0",x"73",x"1B",x"29",x"93",x"01",x"F0",x"59",x"9C",x"0F",x"A9",x"B7",x"04",x"8D",x"1B",x"2B",x"80",x"B0",x"4A",x"5E",x"AD",x"32",x"D8",x"71",x"20",x"14",x"DC",x"D1",x"BC",x"B8",x"4D",x"9F",x"19",x"8F",x"D7",x"3C",x"78",x"AF",x"59",x"12",x"67",x"9A",x"83",x"C9",x"E7",x"C4",x"90",x"0B",x"32",x"88",x"13",x"D8",x"42",x"69",x"A3",x"96",x"69",x"49",x"29",x"49",x"AD",x"6A",x"99",x"AE",x"76",x"CE",x"56",x"89",x"AF",x"64",x"0D",x"4A",x"96",x"6C",x"A9",x"67",x"83",x"6A",x"6B",x"AD",x"67",x"F7",x"86",x"EA",x"22",x"1E",x"A9",x"61",x"A2",x"FC",x"E4",x"8B",x"09",x"30",x"C0",x"BC",x"14",x"DB",x"85",x"04",x"8C",x"B0",x"29",x"B3",x"32",x"65",x"9B",x"9E",x"22",x"AC",x"5C",x"61",x"77",x"CC",x"75",x"62",x"C7",x"5C",x"C3",x"63",x"8A",x"56",x"56",x"64",x"A9",x"39",x"8D",x"65",x"6F",x"29",x"67",x"D0",x"9C",x"96",x"0C",x"F7",x"C9",x"05",x"D9",x"B0",x"20",x"58",x"D3",x"18",x"6D",x"C7",x"99",x"6C",x"65",x"AC",x"C6",x"B9",x"B2",x"61",x"8D",x"29",x"9A",x"68",x"3C",x"69",x"D9",x"B7",x"59",x"97",x"D4",x"45",x"78",x"64",x"A9",x"08",x"9C",x"6B",x"D2",x"CC",x"84",x"DF",x"1F",x"26",x"2F",x"91",x"85",x"37",x"40",x"C0",x"67",x"08",x"C6",x"71",x"38",x"8D",x"E1",x"09",x"1E",x"D0",x"C8",x"C5",x"26",x"F2",x"84",x"34",x"80",x"8F",x"05",x"B2",x"A3",x"71",x"F7",x"6C",x"03",x"A8",x"B1",x"C2",x"E0",x"E9",x"FD",x"E4",x"3A",x"3C",x"D9",x"6D",x"99",x"B0",x"A1",x"11",x"7C",x"A1",x"0D",x"81",x"D1",x"7A",x"6A",x"D4",x"6E",x"8E",x"62",x"D7",x"4C",x"8C",x"08",x"9A",x"64",x"63",x"B0",x"01",x"80",x"F5",x"07",x"95",x"16",x"8F",x"03",x"30",x"3D",x"C7",x"59",x"37",x"EC",x"28",x"80",x"CC",x"65",x"E0",x"91",x"08",x"96",x"80",x"62",x"CE",x"3C",x"49",x"B6",x"04",x"59",x"C2",x"8D",x"8C",x"AB",x"83",x"DB",x"4A",x"03",x"53",x"F8",x"48",x"02",x"98",x"9A",x"24",x"A2",x"07",x"72",x"66",x"AB",x"EC",x"02",x"A3",x"87",x"90",x"50",x"EA",x"BE",x"50",x"B1",x"60",x"08",x"30",x"8B",x"2B",x"D9",x"1A",x"41",x"58",x"8B",x"05",x"7A",x"AE",x"15",x"60",x"EE",x"30",x"ED",x"2C",x"B0",x"4E",x"FC",x"D3",x"12",x"6C",x"08",x"62",x"AA",x"1F",x"FA",x"3B",x"DB",x"98",x"50",x"5F",x"21",x"77",x"34",x"D6",x"A9",x"8F",x"90",x"14",x"57",x"B1",x"BE",x"9C",x"15",x"76",x"90",x"F8",x"FA",x"9C",x"83",x"0C",x"2F",x"41",x"EA",x"84",x"75",x"4E",x"00",x"04",x"34",x"10",x"08",x"F5",x"B9",x"14",x"00",x"28",x"69",x"33",x"67",x"01",x"3A",x"10",x"E3",x"59",x"C9",x"14",x"F0",x"05",x"BF",x"AD",x"08",x"BB",x"2F",x"DE",x"37",x"CF",x"BC",x"2C",x"03",x"40",x"B9",x"A4",x"04",x"06",x"29",x"A9",x"40",x"48",x"83",x"64",x"00",x"78",x"5B",x"67",x"B1",x"E6",x"D3",x"CB",x"58",x"04",x"5C",x"51",x"05",x"24",x"4C",x"DC",x"37",x"ED",x"64",x"C9",x"0D",x"D0",x"1B",x"C8",x"FF",x"04",x"3C",x"BC",x"09",x"F8",x"E4",x"46",x"6D",x"4C",x"F2",x"37",x"77",x"1E",x"02",x"AB",x"D6",x"C6",x"3E",x"71",x"EA",x"C2",x"DA",x"44",x"48",x"24",x"00",x"5E",x"06",x"AB",x"82",x"CD",x"4B",x"80",x"17",x"F4",x"03",x"8A",x"6B",x"69",x"07",x"F8",x"A3",x"DD",x"D4",x"3A",x"EC",x"05",x"5B",x"A8",x"5D",x"A2",x"80",x"8C",x"72",x"9B",x"66",x"D2",x"64",x"2B",x"C6",x"9E",x"71",x"6A",x"A3",x"04",x"88",x"D9",x"B6",x"20",x"D2",x"61",x"70",x"71",x"7B",x"61",x"74",x"92",x"04",x"37",x"5E",x"10",x"D6",x"A0",x"01",x"B9",x"8A",x"8F",x"03",x"62",x"32",x"35",x"F5",x"09",x"4C",x"09",x"74",x"E9",x"B0",x"3C",x"63",x"26",x"E6",x"0B",x"C8",x"4B",x"02",x"CF",x"E1",x"AD",x"0A",x"41",x"FC",x"14",x"D0",x"7A",x"06",x"10",x"3F",x"0C",x"85",x"42",x"C0",x"17",x"A6",x"5F",x"65",x"E5",x"B1",x"1D",x"11",x"C0",x"CF",x"19",x"0B",x"38",x"B7",x"0B",x"F1",x"D3",x"A7",x"80",x"49",x"36",x"E4",x"9D",x"07",x"5B",x"35",x"B5",x"EB",x"CD",x"C3",x"DD",x"80",x"36",x"BB",x"9C",x"C7",x"2D",x"D9",x"87",x"8A",x"09",x"53",x"7B",x"78",x"D4",x"67",x"3C",x"79",x"AE",x"5C",x"3D",x"C5",x"A9",x"20",x"0F",x"F0",x"30",x"74",x"AE",x"6A",x"D0",x"46",x"AA",x"91",x"92",x"56",x"C8",x"D1",x"36",x"B0",x"38",x"35",x"2B",x"10",x"B9",x"CE",x"2C",x"49",x"66",x"52",x"5C",x"CF",x"04",x"3D",x"C5",x"0E",x"89",x"66",x"7D",x"20",x"FF",x"2C",x"A0",x"F8",x"FB",x"B0",x"64",x"9C",x"80",x"C1",x"B8",x"12",x"38",x"D2",x"F1",x"63",x"4E",x"DF",x"2F",x"9C",x"5C",x"33",x"99",x"93",x"31",x"F0",x"2B",x"F8",x"E9",x"75",x"20",x"3B",x"AC",x"76",x"56",x"26",x"7D",x"B1",x"46",x"C2",x"44",x"80",x"C2",x"26",x"29",x"AA",x"D7",x"C8",x"94",x"BA",x"3A",x"CA",x"6B",x"EE",x"2B",x"AD",x"71",x"7D",x"EC",x"8C",x"AC",x"8B",x"56",x"5C",x"4A",x"87",x"6B",x"38",x"0B",x"EF",x"F8",x"07",x"5B",x"70",x"80",x"91",x"04",x"FF",x"12",x"61",x"01",x"0E",x"3A",x"B7",x"C8",x"72",x"22",x"33",x"34",x"14",x"50",x"92",x"EF",x"B6",x"80",x"FE",x"DC",x"90",x"B0",x"37",x"71",x"1B",x"30",x"A3",x"B7",x"99",x"63",x"2F",x"CD",x"16",x"60",x"D7",x"40",x"AD",x"30",x"79",x"79",x"66",x"3E",x"A5",x"40",x"D8",x"A9",x"A0",x"CC",x"0F",x"02",x"7D",x"61",x"F1",x"64",x"63",x"80",x"21",x"F7",x"30",x"87",x"F3",x"03",x"8D",x"43",x"EE",x"D6",x"18",x"58",x"63",x"43",x"55",x"59",x"55",x"21",x"03",x"26",x"D1",x"47",x"EB",x"08",x"07",x"87",x"0F",x"92",x"91",x"B2",x"FA",x"84",x"C8",x"C1",x"30",x"64",x"0C",x"08",x"36",x"41",x"53",x"27",x"B3",x"C5",x"85",x"80",x"87",x"40",x"EF",x"D7",x"F7",x"00",x"57",x"18",x"EB",x"F4",x"13",x"48",x"8A",x"8A",x"1B",x"1C",x"04",x"43",x"21",x"2C",x"96",x"3A",x"81",x"49",x"BC",x"77",x"00",x"5B",x"A9",x"E0",x"C1",x"19",x"2B",x"68",x"C2",x"5B",x"5A",x"BE",x"19",x"71",x"A6",x"8B",x"72",x"72",x"D3",x"1C",x"65",x"FD",x"7D",x"A6",x"54",x"68",x"DF",x"FA",x"8E",x"8E",x"E3",x"F7",x"DC",x"50",x"3A",x"E5",x"0D",x"5A",x"7A",x"29",x"91",x"8D",x"7B",x"5B",x"72",x"7C",x"FA",x"34",x"9A",x"4A",x"9C",x"7E",x"A9",x"01",x"F6",x"88",x"80",x"1B",x"8C",x"30",x"20",x"C4",x"B1",x"C4",x"99",x"CA",x"08",x"8D",x"49",x"CD",x"7E",x"EA",x"01",x"DD",x"F1",x"7F",x"69",x"CD",x"28",x"D0",x"D5",x"D9",x"3E",x"02",x"B9",x"0B",x"D4",x"D0",x"C7",x"9C",x"DB",x"B2",x"10",x"A9",x"0A",x"EA",x"25",x"06",x"D9",x"97",x"10",x"78",x"2D",x"F9",x"29",x"F0",x"D0",x"EA",x"21",x"FC",x"6D",x"92",x"C5",x"8D",x"8A",x"CA",x"61",x"80",x"92",x"76",x"6A",x"98",x"97",x"9A",x"1D",x"F3",x"42",x"BB",x"69",x"38",x"92",x"DC",x"51",x"01",x"90",x"B3",x"46",x"21",x"88",x"88",x"6C",x"03",x"F8",x"60",x"04",x"50",x"C4",x"7D",x"E0",x"FA",x"69",x"07",x"F0",x"33",x"6D",x"1A",x"05",x"2C",x"1E",x"CF",x"4B",x"36",x"65",x"22",x"80",x"92",x"BA",x"2C",x"02",x"6B",x"0E",x"9D",x"4A",x"F0",x"38",x"BF",x"21",x"1E",x"55",x"11",x"F6",x"C7",x"41",x"71",x"1A",x"D8",x"00",x"98",x"11",x"C0",x"14",x"39",x"01",x"13",x"12",x"F8",x"4D",x"90",x"11",x"83",x"DE",x"80",x"C3",x"14",x"3A",x"43",x"3F",x"80",x"3C",x"E0",x"A8",x"18",x"E5",x"21",x"21",x"C8",x"47",x"44",x"F0",x"1A",x"3A",x"E5",x"80",x"32",x"0C",x"80",x"15",x"79",x"8A",x"B8",x"08",x"6D",x"FA",x"68",x"83",x"DC",x"1F",x"34",x"32",x"02",x"13",x"13",x"C8",x"52",x"A6",x"D8",x"52",x"03",x"53",x"10",x"14",x"D8",x"04",x"98",x"84",x"15",x"C0",x"97",x"E2",x"64",x"9E",x"51",x"C0",x"23",x"60",x"1B",x"16",x"4C",x"11",x"10",x"3B",x"6A",x"55",x"82",x"20",x"93",x"DA",x"69",x"A2",x"71",x"FD",x"AF",x"66",x"93",x"AD",x"17",x"38",x"D0",x"3A",x"29",x"5D",x"4A",x"F5",x"B9",x"76",x"47",x"D3",x"D5",x"34",x"A8",x"54",x"E7",x"0B",x"FE",x"40",x"9A",x"F0",x"5C",x"7E",x"C1",x"4E",x"D4",x"84",x"CF",x"9C",x"29",x"7F",x"20",x"43",x"F7",x"62",x"91",x"C1",x"15",x"61",x"6B",x"A2",x"1B",x"4C",x"6E",x"92",x"2B",x"0A",x"05",x"A2",x"CE",x"87",x"94",x"0B",x"2E",x"48",x"88",x"96",x"46",x"03",x"2A",x"04",x"8B",x"F2",x"00",x"3F",x"71",x"07",x"1F",x"60",x"EC",x"DB",x"8D",x"1F",x"CF",x"B0",x"8C",x"67",x"A7",x"23",x"58",x"93",x"AE",x"70",x"35",x"AE",x"4B",x"3B",x"44",x"03",x"90",x"B8",x"2E",x"41",x"14",x"E3",x"94",x"C5",x"A3",x"E1",x"87",x"8B",x"BF",x"71",x"03",x"63",x"02",x"AA",x"D5",x"37",x"50",x"13",x"EE",x"61",x"80",x"6F",x"D1",x"ED",x"98",x"E8",x"3E",x"C7",x"9D",x"56",x"D1",x"08",x"05",x"A3",x"D2",x"04",x"F5",x"E1",x"F4",x"83",x"72",x"67",x"49",x"7A",x"5A",x"66",x"8E",x"76",x"0F",x"64",x"8D",x"8D",x"2E",x"91",x"EA",x"90",x"79",x"8F",x"8E",x"DE",x"16",x"83",x"95",x"7A",x"94",x"49",x"86",x"93",x"9B",x"AD",x"92",x"D2",x"78",x"09",x"D2",x"4F",x"5A",x"09",x"A1",x"41",x"80",x"1F",x"05",x"AE",x"0F",x"02",x"1B",x"B3",x"91",x"3D",x"72",x"F1",x"1A",x"FC",x"E5",x"08",x"00",x"1B",x"67",x"05",x"C7",x"6B",x"EA",x"E7",x"A9",x"02",x"C5",x"49",x"A7",x"E0",x"28",x"67",x"D3",x"AB",x"F3",x"79",x"69",x"71",x"59",x"7D",x"6B",x"E5",x"27",x"B9",x"D7",x"4D",x"75",x"6F",x"2B",x"6F",x"F8",x"AE",x"20",x"BE",x"67",x"60",x"56",x"D2",x"1E",x"6E",x"A9",x"4E",x"45",x"2B",x"EC",x"A9",x"09",x"50",x"68",x"D2",x"8D",x"E2",x"D0",x"B2",x"A4",x"22",x"57",x"2F",x"D6",x"04",x"A0",x"2A",x"FE",x"4A",x"18",x"25",x"BF",x"41",x"FB",x"EB",x"03",x"CE",x"80",x"0B",x"B1",x"41",x"8C",x"9C",x"08",x"B0",x"2E",x"71",x"27",x"A4",x"03",x"F1",x"C2",x"CD",x"5A",x"F4",x"22",x"F1",x"91",x"47",x"3C",x"02",x"CC",x"A9",x"08",x"1F",x"F6",x"2A",x"B0",x"BC",x"03",x"90",x"66",x"48",x"52",x"D2",x"68",x"24",x"CD",x"24",x"64",x"86",x"0B",x"9C",x"2E",x"92",x"0A",x"77",x"9E",x"03",x"8D",x"B0",x"48",x"73",x"70",x"5A",x"82",x"2B",x"4B",x"1C",x"3D",x"D4",x"02",x"8B",x"65",x"96",x"03",x"78",x"FF",x"34",x"26",x"DA",x"08",x"51",x"94",x"D6",x"91",x"11",x"65",x"7E",x"69",x"11",x"22",x"8A",x"18",x"55",x"CE",x"53",x"91",x"F0",x"AB",x"7C",x"38",x"B2",x"DD",x"A9",x"91",x"03",x"47",x"80",x"05",x"5B",x"6C",x"C2",x"3A",x"CE",x"3A",x"BA",x"28",x"D5",x"91",x"29",x"39",x"97",x"FC",x"E1",x"D5",x"91",x"5C",x"A9",x"41",x"F3",x"92",x"05",x"85",x"9E",x"B9",x"F0",x"CD",x"E1",x"9D",x"F2",x"67",x"72",x"43",x"CD",x"35",x"0A",x"6B",x"0C",x"36",x"7E",x"E9",x"BE",x"AA",x"65",x"36",x"54",x"C7",x"94",x"54",x"1D",x"35",x"88",x"D8",x"B8",x"00",x"35",x"54",x"62",x"73",x"63",x"19",x"FC",x"29",x"A9",x"A9",x"01",x"4C",x"B7",x"D9",x"8E",x"B9",x"C3",x"67",x"CC",x"2B",x"5B",x"6D",x"CE",x"9A",x"80",x"0B",x"88",x"E0",x"E4",x"2B",x"E4",x"D0",x"E5",x"9A",x"0D",x"D0",x"0A",x"62",x"10",x"12",x"A3",x"55",x"BB",x"39",x"CC",x"F6",x"26",x"CA",x"42",x"4E",x"10",x"46",x"95",x"81",x"2B",x"B0",x"E7",x"50",x"24",x"09",x"A4",x"42",x"80",x"49",x"95",x"31",x"4F",x"3D",x"4A",x"EB",x"29",x"F9",x"39",x"32",x"A9",x"AB",x"19",x"14",x"A7",x"53",x"90",x"13",x"60",x"7D",x"4D",x"9C",x"FD",x"2C",x"20",x"22",x"63",x"EE",x"2E",x"9E",x"80",x"9E",x"BB",x"DB",x"4E",x"CD",x"BB",x"B0",x"36",x"DA",x"09",x"51",x"A8",x"69",x"42",x"67",x"9F",x"AD",x"9A",x"78",x"5D",x"B7",x"65",x"8E",x"5A",x"8F",x"EF",x"2E",x"B3",x"73",x"3A",x"1D",x"5D",x"80",x"E2",x"C3",x"9A",x"02",x"8B",x"23",x"05",x"90",x"17",x"D7",x"4D",x"39",x"B5",x"36",x"F0",x"B0",x"18",x"71",x"9F",x"3F",x"A3",x"67",x"50",x"4E",x"19",x"0E",x"3E",x"45",x"E9",x"41",x"F0",x"60",x"B4",x"38",x"6E",x"91",x"8E",x"1B",x"97",x"24",x"DC",x"43",x"AD",x"21",x"5E",x"C8",x"A2",x"7C",x"47",x"0F",x"55",x"7C",x"58",x"D5",x"94",x"B1",x"52",x"34",x"78",x"B0",x"27",x"07",x"DB",x"07",x"D0",x"15",x"6B",x"EF",x"78",x"61",x"1F",x"CF",x"67",x"59",x"15",x"0D",x"57",x"11",x"28",x"B7",x"09",x"12",x"80",x"40",x"6C",x"53",x"BF",x"94",x"10",x"93",x"45",x"13",x"43",x"A3",x"4E",x"1E",x"EC",x"49",x"39",x"80",x"23",x"42",x"27",x"29",x"3D",x"40",x"0E",x"38",x"9C",x"D5",x"18",x"A6",x"BA",x"3E",x"87",x"0D",x"6A",x"F3",x"42",x"1C",x"CC",x"42",x"BF",x"02",x"B5",x"CA",x"4C",x"EA",x"CF",x"48",x"0F",x"C5",x"D8",x"51",x"AA",x"8F",x"2E",x"29",x"14",x"55",x"61",x"3E",x"4D",x"57",x"4C",x"6D",x"E4",x"8C",x"92",x"D6",x"69",x"EB",x"E2",x"26",x"85",x"56",x"A8",x"89",x"29",x"8D",x"76",x"78",x"3D",x"A9",x"0F",x"3A",x"3F",x"59",x"9C",x"78",x"20",x"B9",x"20",x"67",x"7E",x"41",x"87",x"CC",x"70",x"AA",x"84",x"24",x"5A",x"BF",x"4B",x"1F",x"3A",x"E0",x"02",x"BF",x"B3",x"B8",x"56",x"45",x"2C",x"CD",x"00",x"B0",x"11",x"4A",x"68",x"43",x"57",x"6C",x"07",x"40",x"6B",x"9C",x"22",x"70",x"0A",x"CD",x"29",x"61",x"D6",x"1C",x"E0",x"2B",x"6C",x"8D",x"77",x"70",x"8A",x"28",x"12",x"9E",x"5F",x"12",x"A4",x"90",x"CB",x"69",x"73",x"AE",x"B6",x"10",x"5B",x"55",x"59",x"18",x"98",x"17",x"EA",x"5B",x"65",x"F0",x"21",x"BC",x"91",x"A9",x"CB",x"18",x"79",x"9E",x"D2",x"11",x"C7",x"2A",x"A2",x"FF",x"86",x"04",x"78",x"2F",x"2E",x"7F",x"DE",x"F8",x"C3",x"2A",x"90",x"D9",x"67",x"5A",x"01",x"4B",x"2E",x"70",x"F0",x"BE",x"61",x"74",x"EB",x"C8",x"55",x"2D",x"10",x"62",x"E0",x"61",x"45",x"4A",x"85",x"92",x"B1",x"59",x"A4",x"62",x"2A",x"FC",x"68",x"D6",x"55",x"7C",x"52",x"6F",x"28",x"5E",x"4C",x"56",x"44",x"BC",x"38",x"DE",x"6E",x"11",x"1A",x"D9",x"20",x"CA",x"0F",x"00",x"B8",x"73",x"30",x"32",x"24",x"77",x"19",x"20",x"AF",x"00",x"8D",x"80",x"D6",x"5D",x"78",x"47",x"40",x"B4",x"25",x"74",x"C9",x"0B",x"B0",x"E6",x"51",x"D3",x"F8",x"18",x"D9",x"A6",x"2F",x"03",x"E0",x"08",x"A9",x"07",x"E5",x"63",x"46",x"4B",x"36",x"0E",x"8D",x"CA",x"33",x"0E",x"48",x"FB",x"73",x"01",x"59",x"3A",x"DD",x"04",x"89",x"6A",x"0E",x"6D",x"6F",x"89",x"C4",x"E5",x"E5",x"F0",x"70",x"D4",x"CE",x"40",x"E2",x"C3",x"92",x"8A",x"E1",x"5E",x"B6",x"BA",x"E5",x"59",x"8A",x"F3",x"58",x"89",x"C1",x"0B",x"85",x"C9",x"08",x"1C",x"7C",x"3F",x"A5",x"02",x"A6",x"03",x"F7",x"28",x"02",x"17",x"3F",x"3B",x"CF",x"2A",x"15",x"94",x"90",x"AC",x"18",x"62",x"FC",x"42",x"A0",x"F7",x"29",x"2A",x"33",x"08",x"28",x"B0",x"63",x"4A",x"1B",x"0E",x"B8",x"0C",x"02",x"2D",x"4C",x"38",x"E9",x"50",x"ED",x"85",x"A9",x"68",x"27",x"2F",x"78",x"22",x"64",x"D1",x"B5",x"D1",x"2C",x"6A",x"CB",x"20",x"92",x"62",x"0C",x"06",x"4F",x"94",x"48",x"A5",x"12",x"05",x"F6",x"18",x"C8",x"0B",x"08",x"B4",x"F1",x"8E",x"2B",x"C8",x"05",x"B1",x"73",x"ED",x"42",x"58",x"1B",x"8A",x"65",x"10",x"A1",x"8D",x"59",x"82",x"8E",x"91",x"42",x"19",x"E4",x"A7",x"1A",x"61",x"4B",x"C1",x"E8",x"B1",x"88",x"A0",x"57",x"4E",x"E6",x"C7",x"67",x"1B",x"21",x"CD",x"DC",x"01",x"9D",x"14",x"87",x"35",x"07",x"D1",x"74",x"12",x"15",x"7C",x"53",x"10",x"BB",x"E3",x"1C",x"E1",x"CC",x"81",x"06",x"1D",x"71",x"1C",x"8A",x"84",x"F8",x"C0",x"80",x"77",x"1E",x"83",x"11",x"04",x"B0",x"A6",x"28",x"32",x"C6",x"1F",x"90",x"02",x"E8",x"BE",x"D4",x"91",x"A8",x"8A",x"7B",x"79",x"AA",x"98",x"F5",x"70",x"2D",x"53",x"0B",x"87",x"07",x"4A",x"E2",x"38",x"6A",x"32",x"0E",x"34",x"70",x"52",x"8B",x"A6",x"A1",x"42",x"3A",x"6A",x"BA",x"6B",x"CD",x"55",x"38",x"CA",x"02",x"EC",x"A1",x"88",x"56",x"B6",x"51",x"5C",x"71",x"5A",x"2A",x"CA",x"69",x"07",x"3B",x"AF",x"8A",x"B5",x"82",x"D9",x"EE",x"A6",x"38",x"33",x"AA",x"6D",x"0A",x"83",x"05",x"2F",x"8A",x"4C",x"FF",x"49",x"DE",x"34",x"14",x"A9",x"47",x"90",x"D1",x"11",x"5B",x"05",x"8A",x"F1",x"35",x"81",x"E0",x"EA",x"A9",x"04",x"28",x"A9",x"2C",x"88",x"81",x"53",x"95",x"54",x"C9",x"4E",x"C6",x"06",x"44",x"63",x"70",x"DE",x"F3",x"F7",x"F0",x"24",x"A6",x"5C",x"1D",x"CC",x"F5",x"66",x"31",x"A3",x"90",x"C4",x"C4",x"F2",x"24",x"C4",x"88",x"5B",x"D0",x"38",x"2E",x"06",x"57",x"05",x"1A",x"B4",x"C7",x"97",x"92",x"61",x"1B",x"B1",x"84",x"D3",x"9F",x"AE",x"A9",x"D2",x"C4",x"66",x"6D",x"52",x"44",x"22",x"EB",x"E7",x"3E",x"10",x"90",x"88",x"5E",x"ED",x"A2",x"6D",x"0B",x"1E",x"B0",x"0A",x"11",x"31",x"1B",x"87",x"A1",x"70",x"53",x"08",x"AE",x"4B",x"09",x"04",x"66",x"4C",x"96",x"87",x"52",x"C6",x"DF",x"2F",x"63",x"A2",x"33",x"38",x"21",x"F2",x"83",x"FA",x"D7",x"69",x"DA",x"34",x"1F",x"5C",x"D3",x"00",x"6C",x"87",x"9D",x"2C",x"0B",x"9C",x"0B",x"80",x"19",x"0B",x"70",x"03",x"0B",x"36",x"E6",x"42",x"02",x"C3",x"65",x"39",x"CE",x"0E",x"00",x"1C",x"36",x"8A",x"35",x"03",x"83",x"AB",x"4C",x"C4",x"4E",x"F4",x"F4",x"65",x"C8",x"F5",x"B8",x"08",x"D0",x"23",x"19",x"54",x"77",x"0C",x"0D",x"83",x"6E",x"00",x"D0",x"A0",x"8B",x"4B",x"71",x"74",x"0F",x"B0",x"EB",x"9E",x"3B",x"F0",x"C8",x"C3",x"32",x"7A",x"A7",x"F8",x"80",x"76",x"C8",x"79",x"32",x"B2",x"02",x"CF",x"E5",x"7C",x"ED",x"64",x"E1",x"74",x"12",x"B7",x"D2",x"5D",x"56",x"96",x"2E",x"A2",x"A1",x"B8",x"07",x"BF",x"66",x"02",x"20",x"37",x"53",x"49",x"3A",x"5D",x"D8",x"A0",x"59",x"B3",x"0D",x"D0",x"03",x"F0",x"BF",x"F9",x"AE",x"E0",x"96",x"65",x"4C",x"7C",x"8B",x"05",x"40",x"68",x"EA",x"78",x"4E",x"31",x"67",x"14",x"68",x"7A",x"4E",x"CB",x"14",x"D9",x"AA",x"89",x"6A",x"D5",x"04",x"B4",x"16",x"4A",x"59",x"8D",x"47",x"D1",x"8E",x"10",x"04",x"BE",x"11",x"95",x"C5",x"CA",x"12",x"64",x"A3",x"85",x"47",x"79",x"F4",x"88",x"4B",x"04",x"7E",x"00",x"B9",x"F4",x"20",x"03",x"87",x"7D",x"3D",x"56",x"BB",x"A0",x"04",x"34",x"AE",x"C1",x"74",x"C9",x"00",x"8A",x"E9",x"7C",x"50",x"A8",x"49",x"80",x"10",x"EB",x"3B",x"8B",x"BB",x"79",x"45",x"12",x"7B",x"C7",x"3D",x"87",x"7B",x"EB",x"18",x"2D",x"D9",x"3D",x"7D",x"C8",x"A7",x"65",x"76",x"0B",x"B2",x"48",x"39",x"5D",x"64",x"D0",x"11",x"0E",x"32",x"61",x"78",x"B8",x"48",x"57",x"6A",x"80",x"B2",x"A0",x"FC",x"CA",x"94",x"50",x"33",x"ED",x"F0",x"7B",x"C4",x"CC",x"B5",x"75",x"00",x"9E",x"A4",x"30",x"18",x"60",x"AA",x"8A",x"02",x"8C",x"A0",x"B0",x"B4",x"AA",x"58",x"8D",x"4B",x"0A",x"6B",x"76",x"D5",x"DD",x"04",x"69",x"C8",x"D3",x"10",x"14",x"9A",x"06",x"1C",x"A3",x"89",x"30",x"0E",x"2D",x"AB",x"CA",x"02",x"29",x"42",x"A9",x"53",x"D0",x"E0",x"4C",x"6D",x"54",x"C0",x"18",x"17",x"09",x"95",x"63",x"6B",x"13",x"01",x"A2",x"DA",x"C8",x"4A",x"74",x"36",x"6A",x"2E",x"EB",x"69",x"5A",x"00",x"EA",x"EB",x"03",x"17",x"DE",x"B4",x"EB",x"01",x"5D",x"58",x"0D",x"38",x"01",x"0D",x"33",x"0D",x"E0",x"06",x"0D",x"08",x"D4",x"42",x"63",x"1A",x"38",x"0B",x"8D",x"A6",x"44",x"68",x"96",x"E6",x"2C",x"74",x"50",x"6A",x"AB",x"01",x"6B",x"66",x"21",x"B0",x"3C",x"57",x"DC",x"41",x"4D",x"B0",x"6D",x"D8",x"E6",x"18",x"0F",x"F9",x"CB",x"A0",x"E6",x"74",x"0E",x"DB",x"30",x"04",x"80",x"0C",x"DC",x"99",x"41",x"91",x"C2",x"AD",x"01",x"3A",x"94",x"00",x"CC",x"EC",x"37",x"87",x"03",x"51",x"09",x"13",x"8B",x"A1",x"A6",x"37",x"4B",x"A5",x"78",x"8E",x"92",x"92",x"B0",x"53",x"E3",x"4C",x"A0",x"4F",x"FD",x"61",x"57",x"A0",x"5E",x"58",x"15",x"06",x"A4",x"62",x"01",x"22",x"16",x"78",x"77",x"26",x"57",x"4E",x"47",x"F1",x"B9",x"60",x"EA",x"81",x"82",x"DE",x"3B",x"15",x"63",x"FF",x"AB",x"20",x"53",x"F3",x"80",x"37",x"07",x"25",x"3D",x"C1",x"F9",x"01",x"BC",x"48",x"1C",x"9C",x"2B",x"AC",x"88",x"92",x"C9",x"6A",x"05",x"7D",x"28",x"E1",x"6E",x"90",x"D9",x"FD",x"0C",x"52",x"5E",x"0C",x"38",x"01",x"0C",x"33",x"0C",x"E0",x"06",x"0C",x"BC",x"DC",x"42",x"26",x"29",x"55",x"91",x"44",x"14",x"C7",x"72",x"64",x"0A",x"65",x"95",x"FF",x"B1",x"0F",x"56",x"37",x"65",x"3A",x"07",x"95",x"95",x"2C",x"13",x"EE",x"81",x"0D",x"02",x"5B",x"78",x"78",x"19",x"09",x"F4",x"80",x"25",x"1A",x"6C",x"C8",x"54",x"1C",x"06",x"AC",x"B6",x"C6",x"8A",x"A6",x"88",x"03",x"34",x"57",x"25",x"8C",x"43",x"E3",x"39",x"7B",x"F7",x"91",x"DE",x"32",x"CB",x"68",x"C1",x"C1",x"E0",x"AE",x"DC",x"CE",x"AB",x"D4",x"D6",x"47",x"8D",x"87",x"67",x"8E",x"88",x"7F",x"E9",x"4C",x"EF",x"50",x"A2",x"96",x"BF",x"98",x"85",x"9A",x"8F",x"80",x"66",x"4F",x"0A",x"BD",x"BA",x"C4",x"9C",x"67",x"59",x"55",x"6A",x"B3",x"AA",x"A2",x"9A",x"56",x"A9",x"65",x"53",x"07",x"9B",x"08",x"50",x"04",x"4F",x"9A",x"17",x"36",x"03",x"4E",x"53",x"0B",x"3D",x"A1",x"4E",x"6C",x"E9",x"A7",x"02",x"86",x"29",x"01",x"0F",x"BB",x"C0",x"0D",x"4C",x"B3",x"B4",x"AD",x"B5",x"65",x"F0",x"FB",x"8D",x"2F",x"9C",x"10",x"D6",x"3B",x"A7",x"1B",x"0E",x"6D",x"60",x"DA",x"40",x"30",x"00",x"C1",x"CE",x"1A",x"01",x"06",x"27",x"86",x"A9",x"B3",x"80",x"8A",x"B2",x"01",x"9C",x"91",x"9D",x"80",x"4E",x"5F",x"BD",x"04",x"1D",x"02",x"67",x"66",x"47",x"8B",x"93",x"65",x"8D",x"BF",x"8E",x"82",x"F6",x"04",x"A5",x"3E",x"1B",x"D5",x"8C",x"56",x"A2",x"74",x"66",x"5D",x"84",x"A9",x"07",x"83",x"92",x"D4",x"03",x"82",x"49",x"64",x"81",x"7D",x"EF",x"39",x"05",x"9A",x"CD",x"60",x"99",x"21",x"05",x"B2",x"5A",x"29",x"A0",x"62",x"41",x"43",x"04",x"B9",x"AF",x"7C",x"90",x"80",x"1F",x"AD",x"E4",x"99",x"15",x"8D",x"CB",x"D5",x"CD",x"12",x"D0",x"F0",x"F9",x"7D",x"90",x"C7",x"D3",x"A9",x"40",x"39",x"87",x"F5",x"C4",x"38",x"B3",x"24",x"78",x"7B",x"41",x"0D",x"E8",x"CF",x"15",x"30",x"5D",x"08",x"4E",x"1E",x"1E",x"A0",x"01",x"AF",x"DC",x"8F",x"14",x"6A",x"61",x"85",x"46",x"D4",x"16",x"CA",x"80",x"70",x"14",x"D6",x"FF",x"49",x"B8",x"8A",x"B9",x"8B",x"EE",x"64",x"34",x"1A",x"67",x"F0",x"EB",x"1C",x"9D",x"8A",x"88",x"A6",x"F9",x"27",x"74",x"5D",x"51",x"01",x"53",x"5A",x"52",x"C1",x"26",x"47",x"4A",x"B4",x"54",x"31",x"61",x"B3",x"5B",x"32",x"4A",x"B2",x"49",x"AD",x"B1",x"78",x"E9",x"AD",x"CE",x"A6",x"65",x"6E",x"66",x"07",x"9D",x"9A",x"17",x"FD",x"31",x"D4",x"10",x"8B",x"27",x"37",x"C5",x"50",x"2D",x"E8",x"03",x"BC",x"0D",x"06",x"53",x"A6",x"07",x"D2",x"C9",x"92",x"64",x"8A",x"04",x"97",x"C3",x"70",x"E9",x"00",x"DD",x"B0",x"3B",x"93",x"75",x"08",x"91",x"A3",x"78",x"2C",x"DF",x"0C",x"65",x"F4",x"16",x"27",x"35",x"C7",x"80",x"04",x"A9",x"22",x"A2",x"76",x"7E",x"A3",x"D0",x"49",x"97",x"82",x"33",x"D6",x"0D",x"C1",x"B5",x"7C",x"83",x"2C",x"5E",x"AF",x"D0",x"82",x"74",x"B6",x"60",x"96",x"21",x"AD",x"24",x"67",x"04",x"2F",x"88",x"C4",x"80",x"8B",x"48",x"61",x"72",x"9C",x"18",x"1A",x"D0",x"4E",x"51",x"8A",x"88",x"5A",x"02",x"43",x"15",x"03",x"6B",x"A5",x"04",x"AB",x"AD",x"7B",x"C8",x"AE",x"7C",x"D2",x"75",x"18",x"B3",x"E7",x"C8",x"6C",x"A7",x"BC",x"7A",x"65",x"A5",x"76",x"78",x"B9",x"20",x"3F",x"6A",x"4C",x"F8",x"55",x"FC",x"0D",x"43",x"9D",x"51",x"00",x"F0",x"8A",x"1C",x"EC",x"1C",x"AA",x"02",x"38",x"07",x"21",x"15",x"09",x"AA",x"AD",x"92",x"0A",x"A2",x"C3",x"A9",x"FB",x"50",x"47",x"80",x"8A",x"3D",x"AD",x"AE",x"DF",x"CD",x"38",x"E9",x"8E",x"B0",x"01",x"CA",x"8D",x"FE",x"8E",x"8E",x"AD",x"85",x"2D",x"0D",x"86",x"7D",x"D0",x"7D",x"A6",x"03",x"56",x"FB",x"85",x"40",x"D0",x"E0",x"E8",x"71",x"C9",x"01",x"F0",x"6A",x"F8",x"07",x"03",x"D0",x"C1",x"B3",x"7A",x"AB",x"0B",x"B0",x"79",x"B5",x"B3",x"B2",x"0A",x"29",x"E8",x"67",x"D0",x"2C",x"20",x"49",x"63",x"7F",x"78",x"15",x"05",x"B6",x"77",x"85",x"D6",x"AE",x"76",x"D6",x"AD",x"A1",x"75",x"A0",x"64",x"20",x"7D",x"6A",x"A9",x"91",x"FB",x"4E",x"79",x"04",x"A3",x"64",x"05",x"B3",x"7B",x"6A",x"A2",x"FF",x"BE",x"2E",x"71",x"2D",x"D5",x"80",x"1E",x"AD",x"1F",x"1A",x"29",x"0F",x"8D",x"FB",x"D0",x"20",x"68",x"4A",x"51",x"C3",x"D1",x"DC",x"A0",x"04",x"B1",x"02",x"F2",x"CA",x"36",x"03",x"49",x"E1",x"54",x"14",x"4D",x"4E",x"0A",x"56",x"0C",x"30",x"CA",x"AA",x"6A",x"54",x"82",x"CB",x"2A",x"89",x"BA",x"07",x"D8",x"5A",x"20",x"28",x"07",x"E3",x"63",x"7C",x"4B",x"7B",x"CE",x"EE",x"EC",x"74",x"54",x"42",x"02",x"28",x"C7",x"49",x"B7",x"09",x"20",x"21",x"6C",x"58",x"5F",x"78",x"97",x"07",x"84",x"76",x"34",x"0F",x"A0",x"E0",x"25",x"14",x"08",x"34",x"F0",x"A0",x"E0",x"D7",x"FF",x"4A",x"84",x"1D",x"30",x"22",x"28",x"53",x"20",x"E0",x"E8",x"62",x"38",x"78",x"A3",x"48",x"58",x"D8",x"C0",x"FF",x"B7",x"29",x"66",x"76",x"F4",x"CF",x"E4",x"AA",x"29",x"6A",x"F8",x"E0",x"7D",x"DC",x"55",x"53",x"FC",x"7C",x"1C",x"04",x"F4",x"87",x"9B",x"22",x"A8",x"70",x"69",x"C3",x"01",x"26",x"6C",x"B0",x"4F",x"99",x"1C",x"22",x"58",x"44",x"F0",x"34",x"88",x"70",x"27",x"88",x"90",x"40",x"47",x"13",x"54",x"55",x"BA",x"1D",x"52",x"5E",x"A5",x"8A",x"00",x"27",x"8E",x"0A",x"25",x"95",x"0C",x"08",x"30",x"9D",x"47",x"83",x"B3",x"3F",x"E8",x"97",x"C5",x"43",x"A8",x"B7",x"B9",x"28",x"47",x"D9",x"95",x"CC",x"C6",x"A0",x"A8",x"FE",x"29",x"37",x"84",x"AB",x"C5",x"C7",x"CC",x"10",x"DF",x"9C",x"A3",x"A6",x"05",x"92",x"04",x"FE",x"48",x"C8",x"6E",x"7C",x"A5",x"B7",x"24",x"F8",x"C4",x"E7",x"EF",x"CE",x"8C",x"E8",x"2B",x"78",x"70",x"CE",x"CC",x"7E",x"F9",x"06",x"F5",x"6F",x"32",x"C4",x"42",x"20",x"EF",x"A6",x"9A",x"8C",x"28",x"27",x"33",x"85",x"FE",x"72",x"93",x"10",x"92",x"32",x"10",x"60",x"47",x"6F",x"05",x"C0",x"D8",x"65",x"04",x"66",x"93",x"93",x"80",x"FD",x"36",x"FC",x"EC",x"7F",x"33",x"70",x"81",x"E6",x"40",x"38",x"60",x"7C",x"9D",x"FC",x"9A",x"9F",x"A1",x"1C",x"3C",x"CC",x"FE",x"7E",x"EC",x"33",x"CC",x"0C",x"A0",x"8C",x"4F",x"7D",x"26",x"CF",x"57",x"6B",x"89",x"13",x"8E",x"60",x"AE",x"4D",x"B2",x"A5",x"F2",x"C0",x"39",x"14",x"27",x"13",x"23",x"62",x"64",x"30",x"14",x"CE",x"0C",x"13",x"2C",x"8D",x"C3",x"59",x"64",x"98",x"83",x"58",x"50",x"32",x"3F",x"53",x"E3",x"34",x"FD",x"A4",x"F8",x"3F",x"A1",x"1A",x"AF",x"7A",x"E9",x"0C",x"C9",x"C1",x"88",x"4E",x"83",x"3F",x"B4",x"A8",x"12",x"78",x"3F",x"15",x"3C",x"81",x"D7",x"CD",x"70",x"E8",x"69",x"13",x"B0",x"BB",x"35",x"C0",x"46",x"F8",x"80",x"3F",x"7A",x"50",x"9D",x"FD",x"92",x"06",x"50",x"87",x"D1",x"F1",x"B9",x"CF",x"3F",x"B4",x"80",x"EC",x"64",x"18",x"D3",x"CC",x"C0",x"0C",x"C5",x"E0",x"3F",x"52",x"0B",x"80",x"B5",x"45",x"46",x"0C",x"3F",x"D5",x"B3",x"60",x"3C",x"FF",x"C0",x"C1",x"60",x"11",x"B7",x"20",x"37",x"C3",x"C5",x"8F",x"7C",x"E2",x"63",x"80",x"3D",x"26",x"6E",x"26",x"53",x"6F",x"86",x"1D",x"0E",x"23",x"D6",x"7A",x"F3",x"CA",x"98",x"4E",x"C4",x"67",x"6E",x"49",x"C9",x"9C",x"48",x"DF",x"80",x"E1",x"CD",x"33",x"B6",x"45",x"78",x"6C",x"9F",x"38",x"90",x"C6",x"9C",x"93",x"71",x"7F",x"6B",x"0D",x"63",x"FA",x"28",x"C6",x"CA",x"77",x"30",x"41",x"2A",x"7C",x"D6",x"31",x"12",x"8C",x"06",x"54",x"38",x"08",x"0B",x"3D",x"30",x"35",x"3E",x"6F",x"BD",x"06",x"CF",x"5D",x"09",x"7E",x"65",x"22",x"0E",x"0F",x"85",x"6B",x"27",x"45",x"67",x"07",x"63",x"6B",x"7F",x"3E",x"36",x"F9",x"87",x"89",x"18",x"3C",x"9E",x"76",x"5F",x"04",x"1B",x"D5",x"44",x"35",x"D7",x"7E",x"B6",x"44",x"86",x"21",x"03",x"82",x"88",x"D2",x"AA",x"04",x"0C",x"0B",x"E1",x"95",x"93",x"32",x"74",x"2C",x"BE",x"03",x"58",x"01",x"82",x"FE",x"F6",x"41",x"40",x"DC",x"4F",x"E4",x"31",x"47",x"F3",x"18",x"66",x"F3",x"6B",x"50",x"7B",x"11",x"69",x"F3",x"33",x"07",x"62",x"7A",x"99",x"5F",x"F7",x"6A",x"AA",x"5B",x"87",x"44",x"7C",x"1E",x"1B",x"8A",x"48",x"6E",x"19",x"D1",x"37",x"01",x"0C",x"65",x"92",x"13",x"89",x"F0",x"D8",x"3E",x"11",x"80",x"C0",x"C9",x"DA",x"A3",x"EE",x"05",x"69",x"D6",x"A1",x"57",x"23",x"D3",x"DC",x"8A",x"3D",x"8F",x"08",x"B0",x"1D",x"2D",x"AF",x"54",x"14",x"D4",x"D8",x"6C",x"2F",x"72",x"35",x"F8",x"47",x"44",x"B3",x"C0",x"E0",x"78",x"3B",x"1C",x"F8",x"F4",x"DB",x"00",x"F3",x"D9",x"61",x"58",x"E6",x"B3",x"58",x"6B",x"22",x"69",x"4B",x"D6",x"42",x"FE",x"EE",x"C6",x"3F",x"08",x"66",x"2C",x"61",x"59",x"2A",x"DC",x"78",x"3F",x"0D",x"81",x"18",x"30",x"77",x"EC",x"7D",x"08",x"60",x"58",x"D1",x"11",x"A1",x"02",x"18",x"98",x"1F",x"2A",x"7C",x"A1",x"00",x"79",x"E0",x"44",x"FE",x"7E",x"20",x"07",x"14",x"5C",x"38",x"C0",x"AA",x"3A",x"44",x"C9",x"48",x"C9",x"6C",x"40",x"BF",x"68",x"F0",x"42",x"60",x"FC",x"8F",x"49",x"24",x"5A",x"D0",x"2B",x"82",x"44",x"6C",x"F2",x"96",x"1B",x"18",x"6F",x"18",x"9C",x"64",x"90",x"83",x"98",x"D9",x"92",x"AB",x"36",x"37",x"A2",x"B2",x"C6",x"37",x"02",x"67",x"08",x"A3",x"38",x"A6",x"8E",x"99",x"A2",x"6E",x"62",x"30",x"7C",x"04",x"2B",x"60",x"1A",x"45",x"35",x"41",x"B2",x"AA",x"44",x"17",x"38",x"90",x"80",x"79",x"55",x"10",x"36",x"41",x"6D",x"3A",x"40",x"E5",x"61",x"02",x"D2",x"B6",x"82",x"08",x"89",x"72",x"64",x"38",x"24",x"B6",x"CB",x"7C",x"42",x"E8",x"68",x"03",x"28",x"F6",x"40",x"00",x"0A",x"C2",x"18",x"04",x"FD",x"42",x"09",x"60",x"05",x"B6",x"B7",x"31",x"09",x"62",x"30",x"0A",x"98",x"C2",x"45",x"12",x"24",x"4F",x"87",x"26",x"A9",x"0F",x"42",x"C4",x"48",x"56",x"22",x"F9",x"86",x"A3",x"C2",x"AD",x"44",x"C8",x"52",x"E6",x"4A",x"84",x"7F",x"B0",x"36",x"60",x"DB",x"24",x"4F",x"72",x"28",x"2E",x"BB",x"43",x"01",x"E4",x"1D",x"64",x"8A",x"98",x"1F",x"48",x"8A",x"08",x"A2",x"0C",x"30",x"94",x"21",x"FC",x"CC",x"37",x"3E",x"85",x"28",x"4E",x"9E",x"88",x"8E",x"6E",x"4D",x"C0",x"35",x"D4",x"89",x"40",x"BE",x"76",x"30",x"5E",x"3B",x"14",x"AF",x"1D",x"0A",x"D4",x"02",x"60",x"7C",x"F2",x"DB",x"0E",x"C6",x"DB",x"0E",x"85",x"64",x"28",x"82",x"58",x"3C",x"13",x"68",x"EC",x"64",x"A1",x"F8",x"7D",x"11",x"4A",x"68",x"58",x"48",x"FA",x"DD",x"0E",x"C6",x"E3",x"0E",x"C5",x"6A",x"87",x"28",x"50",x"E2",x"43",x"D1",x"D9",x"04",x"AC",x"6E",x"D7",x"64",x"8A",x"56",x"44",x"F6",x"A7",x"1A",x"95",x"2C",x"34",x"24",x"58",x"FE",x"48",x"0E",x"20",x"8C",x"8F",x"E2",x"87",x"C5",x"D3",x"00",x"CC",x"78",x"E4",x"0F",x"6C",x"38",x"CE",x"D7",x"84",x"F8",x"14",x"CC",x"FC",x"1A",x"C0",x"34",x"6D",x"02",x"81",x"64",x"68",x"06",x"26",x"20",x"8D",x"10",x"8B",x"07",x"E3",x"E7",x"0C",x"EA",x"48",x"79",x"30",x"F2",x"78",x"08",x"76",x"CC",x"7C",x"F4",x"29",x"EC",x"32",x"39",x"90",x"F4",x"D4",x"4D",x"C0",x"32",x"13",x"20",x"7D",x"25",x"87",x"02",x"6C",x"8F",x"02",x"6C",x"78",x"2B",x"BB",x"55",x"7E",x"60",x"3C",x"FC",x"20",x"1E",x"0C",x"B7",x"1D",x"0A",x"E9",x"50",x"F8",x"CD",x"33",x"60",x"AA",x"45",x"20",x"50",x"4B",x"24",x"18",x"D0",x"2F",x"7C",x"A6",x"8D",x"7C",x"C6",x"3A",x"14",x"6F",x"5B",x"10",x"3C",x"18",x"14",x"28",x"1B",x"66",x"3A",x"25",x"93",x"11",x"3C",x"59",x"36",x"20",x"7C",x"53",x"03",x"56",x"3A",x"4C",x"54",x"64",x"B8",x"FD",x"D7",x"0E",x"20",x"8C",x"AC",x"43",x"10",x"28",x"F1",x"41",x"44",x"B1",x"02",x"C6",x"7E",x"C8",x"08",x"AE",x"10",x"1F",x"05",x"8B",x"92",x"48",x"A0",x"70",x"40",x"87",x"24",x"EA",x"BA",x"3E",x"0C",x"CF",x"78",x"45",x"C4",x"20",x"8F",x"DE",x"21",x"AA",x"97",x"F0",x"E3",x"3A",x"BC",x"69",x"C5",x"B3",x"FF",x"9D",x"D4",x"BF",x"36",x"CE",x"54",x"D0",x"FD",x"28",x"61",x"2B",x"B5",x"8D",x"AD",x"C8",x"7E",x"A9",x"90",x"DD",x"A2",x"E3",x"20",x"9B",x"5E",x"EF",x"33",x"A5",x"A9",x"16",x"78",x"33",x"5C",x"17",x"60",x"3E",x"11",x"15",x"9C",x"62",x"AD",x"73",x"6A",x"AF",x"CD",x"6B",x"E7",x"96",x"62",x"7C",x"4E",x"E1",x"C9",x"20",x"45",x"5E",x"67",x"F3",x"2C",x"0D",x"13",x"4D",x"16",x"AD",x"D2",x"0A",x"84",x"0B",x"F3",x"D1",x"4A",x"EE",x"30",x"90",x"2C",x"EF",x"C9",x"9B",x"B0",x"46",x"70",x"24",x"48",x"67",x"66",x"30",x"8C",x"69",x"C2",x"0C",x"B8",x"B8",x"27",x"A6",x"7B",x"68",x"65",x"8E",x"60",x"90",x"D1",x"DD",x"E6",x"B0",x"AB",x"CD",x"9A",x"6B",x"AC",x"44",x"3A",x"49",x"99",x"CD",x"89",x"60",x"A9",x"9D",x"7A",x"9F",x"18",x"6D",x"B7",x"9C",x"E9",x"87",x"C5",x"20",x"85",x"A6",x"1B",x"DD",x"4C",x"53",x"A3",x"D5",x"5E",x"96",x"56",x"F8",x"B1",x"EE",x"17",x"BC",x"F3",x"D1",x"FF",x"D0",x"5E",x"B1",x"6E",x"35",x"08",x"B0",x"AE",x"50",x"5C",x"FF",x"DF",x"4C",x"92",x"B3",x"8E",x"61",x"41",x"67",x"84",x"78",x"4B",x"4F",x"66",x"20",x"C2",x"5E",x"FA",x"8D",x"4C",x"82",x"67",x"EE",x"48",x"6D",x"B9",x"DA",x"00",x"99",x"D7",x"9B",x"2E",x"EE",x"F7",x"68",x"EF",x"16",x"5A",x"17",x"18",x"4F",x"19",x"A6",x"3B",x"F6",x"B0",x"86",x"1B",x"D7",x"1E",x"97",x"91",x"52",x"3A",x"32",x"AB",x"66",x"8D",x"33",x"CA",x"79",x"27",x"95",x"0A",x"1D",x"85",x"B3",x"B9",x"34",x"18",x"47",x"0B",x"53",x"A9",x"2E",x"DC",x"F5",x"DC",x"1C",x"EC",x"98",x"DB",x"65",x"1A",x"18",x"BD",x"55",x"15",x"38",x"A6",x"0A",x"B5",x"6A",x"A5",x"19",x"E5",x"0B",x"85",x"0D",x"FD",x"0C",x"AD",x"F0",x"25",x"20",x"2F",x"63",x"23",x"FF",x"AF",x"1B",x"1A",x"9E",x"0B",x"E7",x"0A",x"49",x"30",x"0D",x"FF",x"69",x"0C",x"26",x"D3",x"27",x"31",x"E5",x"EA",x"24",x"5E",x"AA",x"FB",x"61",x"A2",x"05",x"BD",x"8A",x"F7",x"7F",x"95",x"16",x"6F",x"F8",x"60",x"ED",x"C2",x"A0",x"25",x"90",x"AF",x"14",x"32",x"43",x"75",x"F3",x"6E",x"0B",x"9D",x"79",x"CA",x"B3",x"10",x"FA",x"D3",x"22",x"2D",x"91",x"CB",x"19",x"5B",x"2B",x"92",x"CB",x"10",x"5B",x"20",x"05",x"AB",x"CB",x"3D",x"07",x"B2",x"23",x"AE",x"E6",x"45",x"81",x"36",x"CF",x"5F",x"C7",x"C9",x"BA",x"30",x"E7",x"55",x"72",x"8E",x"88",x"95",x"7F",x"37",x"18",x"4C",x"96",x"34",x"97",x"B3",x"C2",x"8C",x"2E",x"0C",x"2E",x"62",x"1B",x"45",x"C8",x"09",x"2A",x"69",x"DF",x"01",x"C9",x"29",x"4C",x"3F",x"60",x"79",x"7A",x"0D",x"DC",x"8E",x"FD",x"75",x"B1",x"18",x"5A",x"D7",x"19",x"5A",x"48",x"15",x"6B",x"54",x"11",x"AD",x"4A",x"75",x"08",x"B4",x"CC",x"12",x"4C",x"91",x"0B",x"0F",x"55",x"9C",x"9A",x"14",x"4C",x"99",x"45",x"C9",x"DD",x"9C",x"9D",x"5E",x"AA",x"57",x"A2",x"BB",x"DE",x"28",x"54",x"56",x"43",x"0E",x"AD",x"DB",x"9D",x"99",x"87",x"34",x"9E",x"B3",x"43",x"44",x"44",x"4F",x"49",x"D0",x"2D",x"5E",x"00",x"93",x"AB",x"61",x"20",x"AD",x"92",x"0E",x"02",x"A2",x"DA",x"2B",x"8E",x"67",x"66",x"24",x"A4",x"05",x"30",x"0B",x"AC",x"9B",x"FF",x"28",x"8C",x"9D",x"59",x"EE",x"9C",x"7F",x"7A",x"0A",x"1D",x"C5",x"4E",x"58",x"15",x"69",x"34",x"49",x"36",x"08",x"C9",x"F2",x"1A",x"F2",x"AD",x"CF",x"39",x"C9",x"4F",x"F9",x"6E",x"20",x"5C",x"5E",x"AC",x"CF",x"4B",x"17",x"48",x"73",x"A6",x"0F",x"09",x"39",x"06",x"C5",x"55",x"68",x"88",x"40",x"7E",x"20",x"FD",x"5E",x"87",x"50",x"99",x"D0",x"65",x"C1",x"A5",x"9A",x"4E",x"E8",x"8E",x"BB",x"A9",x"D9",x"C1",x"27",x"C9",x"53",x"E6",x"DD",x"20",x"6E",x"5E",x"EF",x"8D",x"8E",x"2F",x"DF",x"1C",x"55",x"D0",x"0B",x"73",x"99",x"89",x"64",x"04",x"48",x"C0",x"C2",x"E6",x"C9",x"D8",x"D0",x"29",x"48",x"FB",x"AD",x"94",x"F3",x"0A",x"D9",x"30",x"4A",x"A9",x"90",x"D8",x"B8",x"AB",x"44",x"51",x"5E",x"A0",x"20",x"DD",x"0A",x"5F",x"68",x"C9",x"F7",x"58",x"16",x"7D",x"0E",x"41",x"6B",x"63",x"69",x"61",x"E9",x"5F",x"AD",x"B1",x"B2",x"AE",x"B2",x"F4",x"B1",x"2B",x"6B",x"8D",x"77",x"D0",x"8E",x"B4",x"EE",x"AC",x"0D",x"58",x"CD",x"F0",x"15",x"AE",x"98",x"5E",x"EC",x"74",x"AD",x"B3",x"99",x"47",x"A8",x"4B",x"06",x"8E",x"E6",x"8C",x"8C",x"ED",x"38",x"D8",x"96",x"4A",x"B3",x"EC",x"AA",x"AD",x"34",x"67",x"ED",x"B4",x"BF",x"E0",x"56",x"30",x"BC",x"97",x"B2",x"AB",x"C2",x"8D",x"96",x"B2",x"54",x"D0",x"2A",x"A6",x"E5",x"B6",x"AD",x"91",x"7F",x"5B",x"EE",x"20",x"DA",x"5E",x"4C",x"4A",x"FB",x"5F",x"B5",x"2B",x"BD",x"05",x"2E",x"B6",x"7F",x"6B",x"50",x"E4",x"D4",x"18",x"E1",x"2B",x"69",x"F4",x"C5",x"77",x"F0",x"16",x"ED",x"41",x"67",x"79",x"18",x"BE",x"98",x"65",x"EB",x"70",x"4F",x"94",x"68",x"54",x"4C",x"C3",x"00",x"C8",x"08",x"0A",x"07",x"59",x"1C",x"44",x"0E",x"52",x"0E",x"43",x"41",x"C3",x"FD",x"A8",x"19",x"0A",x"23",x"58",x"57",x"FD",x"9E",x"BA",x"5A",x"70",x"A6",x"5B",x"F5",x"0D",x"B4",x"E8",x"F4",x"44",x"11",x"FF",x"9B",x"8B",x"7F",x"B0",x"02",x"16",x"6B",x"01",x"34",x"06",x"AA",x"AD",x"2B",x"FD",x"91",x"A7",x"34",x"35",x"5E",x"C4",x"AD",x"36",x"2C",x"AE",x"37",x"79",x"BD",x"86",x"63",x"E6",x"FF",x"19",x"5D",x"00",x"49",x"CB",x"77",x"08",x"DA",x"3E",x"36",x"24",x"15",x"59",x"9C",x"6F",x"76",x"90",x"05",x"3D",x"40",x"4A",x"18",x"29",x"0F",x"FE",x"55",x"64",x"A2",x"69",x"38",x"57",x"D3",x"36",x"A4",x"C5",x"28",x"BB",x"F4",x"30",x"88",x"88",x"71",x"60",x"3D",x"04",x"7C",x"05",x"F8",x"06",x"F0",x"07",x"21",x"E3",x"74",x"A0",x"FB",x"C7",x"02",x"ED",x"D8",x"73",x"24",x"5B",x"5A",x"18",x"BD",x"5D",x"EE",x"79",x"79",x"E8",x"BB",x"E0",x"08",x"90",x"F6",x"60",x"8C",x"FF",x"28",x"D8",x"AD",x"92",x"2E",x"18",x"52",x"6B",x"4B",x"68",x"90",x"AC",x"01",x"E8",x"03",x"97",x"AF",x"19",x"AD",x"10",x"F9",x"31",x"8C",x"49",x"89",x"6C",x"AC",x"B7",x"AF",x"5A",x"8D",x"91",x"8E",x"E7",x"86",x"C5",x"45",x"29",x"01",x"6C",x"E9",x"A9",x"10",x"20",x"C9",x"61",x"AA",x"FE",x"5F",x"52",x"29",x"2C",x"94",x"F1",x"5E",x"6D",x"3D",x"25",x"57",x"6A",x"5E",x"62",x"9A",x"76",x"51",x"09",x"97",x"95",x"68",x"E0",x"E6",x"C3",x"0E",x"C9",x"00",x"D0",x"9E",x"B5",x"43",x"0A",x"54",x"6E",x"20",x"72",x"6C",x"72",x"79",x"18",x"C9",x"CA",x"7E",x"14",x"B6",x"B8",x"55",x"CC",x"AD",x"B9",x"7F",x"C3",x"75",x"3F",x"C6",x"09",x"2B",x"DD",x"D0",x"95",x"A5",x"7D",x"A9",x"69",x"5F",x"8E",x"C1",x"65",x"20",x"C4",x"6B",x"7E",x"7B",x"5B",x"3E",x"6F",x"DD",x"8E",x"CC",x"F9",x"C8",x"A1",x"C8",x"19",x"95",x"09",x"E2",x"B0",x"80",x"BC",x"F3",x"69",x"5A",x"B2",x"FD",x"52",x"8B",x"73",x"42",x"D0",x"96",x"0C",x"16",x"8F",x"01",x"05",x"79",x"F0",x"C5",x"A2",x"18",x"4F",x"5A",x"A2",x"04",x"9C",x"05",x"E7",x"06",x"79",x"07",x"12",x"36",x"E6",x"4F",x"62",x"94",x"5A",x"81",x"33",x"D3",x"88",x"CA",x"95",x"D1",x"53",x"4C",x"3B",x"69",x"54",x"18",x"6B",x"A1",x"12",x"0E",x"23",x"33",x"88",x"91",x"29",x"6D",x"22",x"75",x"18",x"6F",x"54",x"E3",x"30",x"34",x"83",x"20",x"64",x"57",x"46",x"07",x"91",x"E3",x"C0",x"02",x"B3",x"1B",x"7B",x"C3",x"33",x"AA",x"2C",x"D9",x"44",x"66",x"4F",x"A9",x"46",x"31",x"AD",x"6D",x"09",x"46",x"86",x"78",x"C4",x"4C",x"A2",x"D0",x"03",x"C5",x"40",x"8A",x"36",x"24",x"26",x"6C",x"CD",x"4D",x"05",x"5B",x"22",x"04",x"CF",x"0C",x"6A",x"0B",x"98",x"D0",x"4B",x"C5",x"0A",x"CD",x"24",x"F0",x"88",x"B0",x"AF",x"03",x"A5",x"96",x"69",x"B4",x"50",x"A4",x"04",x"09",x"C9",x"08",x"20",x"D6",x"BF",x"28",x"B5",x"37",x"78",x"72",x"0A",x"D3",x"72",x"CD",x"05",x"49",x"90",x"D0",x"86",x"88",x"AA",x"AD",x"E3",x"E1",x"67",x"14",x"20",x"38",x"93",x"DA",x"B0",x"0D",x"DE",x"CA",x"E0",x"FF",x"08",x"AF",x"55",x"E4",x"68",x"C6",x"69",x"D7",x"9A",x"6F",x"68",x"CE",x"84",x"A5",x"C5",x"D0",x"F9",x"09",x"E8",x"06",x"AE",x"93",x"AB",x"9F",x"C2",x"1A",x"A1",x"D1",x"CF",x"59",x"51",x"0E",x"C5",x"0F",x"92",x"60",x"10",x"54",x"EA",x"95",x"F8",x"59",x"94",x"68",x"91",x"8D",x"35",x"3B",x"46",x"15",x"EF",x"14",x"50",x"13",x"6A",x"E9",x"68",x"BC",x"0B",x"66",x"0A",x"90",x"17",x"F9",x"18",x"0E",x"A9",x"48",x"0F",x"6B",x"15",x"13",x"D5",x"10",x"5A",x"45",x"C4",x"DE",x"11",x"65",x"EB",x"08",x"D8",x"3B",x"10",x"B9",x"D5",x"F7",x"89",x"18",x"58",x"20",x"01",x"A1",x"1B",x"C6",x"32",x"2C",x"87",x"21",x"AD",x"6D",x"88",x"69",x"00",x"EE",x"00",x"4E",x"D8",x"05",x"4A",x"CA",x"9D",x"33",x"A2",x"6D",x"4C",x"5A",x"64",x"FF",x"71",x"2C",x"B1",x"48",x"8A",x"20",x"15",x"63",x"7F",x"5F",x"05",x"92",x"20",x"6A",x"78",x"6B",x"A8",x"3D",x"85",x"06",x"86",x"07",x"7E",x"8A",x"08",x"A4",x"DB",x"28",x"27",x"60",x"5A",x"09",x"2B",x"95",x"08",x"D4",x"A6",x"07",x"DB",x"A5",x"06",x"60",x"29",x"1F",x"BF",x"3C",x"31",x"D2",x"D5",x"D8",x"F0",x"0E",x"A8",x"BD",x"08",x"88",x"E3",x"77",x"C4",x"68",x"E8",x"14",x"2C",x"9E",x"A2",x"96",x"71",x"CB",x"10",x"12",x"38",x"01",x"9A",x"76",x"5E",x"54",x"4D",x"84",x"0B",x"C6",x"91",x"B1",x"21",x"C3",x"66",x"A5",x"45",x"A2",x"62",x"AA",x"11",x"33",x"61",x"66",x"33",x"53",x"0A",x"69",x"33",x"B4",x"D8",x"00",x"62",x"26",x"D7",x"06",x"15",x"E5",x"B7",x"57",x"4E",x"BB",x"6E",x"9D",x"CF",x"2F",x"12",x"B0",x"C9",x"0D",x"A8",x"98",x"36",x"DF",x"F9",x"DB",x"CF",x"62",x"87",x"BB",x"29",x"A5",x"BC",x"EC",x"04",x"86",x"5C",x"60",x"0A",x"8A",x"A6",x"74",x"D6",x"B9",x"C0",x"2D",x"39",x"B6",x"04",x"E2",x"22",x"0A",x"11",x"A7",x"E0",x"80",x"AD",x"FF",x"A0",x"0B",x"ED",x"58",x"76",x"DA",x"63",x"88",x"F8",x"AB",x"4C",x"B9",x"67",x"8A",x"10",x"1D",x"A9",x"2D",x"FF",x"84",x"2B",x"5C",x"0C",x"5E",x"CD",x"0D",x"64",x"AD",x"79",x"13",x"66",x"8D",x"CD",x"4C",x"85",x"99",x"70",x"29",x"67",x"0B",x"48",x"2B",x"E8",x"70",x"0E",x"1A",x"C5",x"C2",x"A9",x"12",x"AD",x"C4",x"EC",x"A8",x"B9",x"F3",x"76",x"48",x"68",x"B2",x"0B",x"D5",x"04",x"50",x"05",x"D0",x"D9",x"A7",x"9E",x"6D",x"F9",x"03",x"DF",x"AE",x"F8",x"3C",x"DB",x"4C",x"44",x"47",x"43",x"80",x"A7",x"0E",x"86",x"FA",x"CF",x"04",x"4E",x"4F",x"58",x"B8",x"BB",x"63",x"0E",x"6B",x"C0",x"2B",x"0B",x"09",x"04",x"B1",x"26",x"96",x"41",x"67",x"48",x"A9",x"F2",x"E2",x"16",x"CD",x"A0",x"20",x"C8",x"1F",x"78",x"42",x"04",x"05",x"A5",x"2A",x"23",x"57",x"14",x"68",x"15",x"A7",x"F5",x"0E",x"76",x"64",x"4A",x"06",x"71",x"0F",x"58",x"00",x"15",x"8A",x"37",x"0E",x"A9",x"A7",x"9B",x"4A",x"0F",x"BD",x"3C",x"B9",x"94",x"F9",x"5B",x"F9",x"03",x"30",x"91",x"DC",x"0C",x"60",x"7D",x"90",x"26",x"8E",x"26",x"86",x"56",x"20",x"1D",x"65",x"4C",x"5F",x"EF",x"A5",x"76",x"04",x"84",x"D1",x"05",x"CF",x"AB",x"20",x"F3",x"67",x"F4",x"14",x"5A",x"04",x"47",x"15",x"42",x"FD",x"3E",x"96",x"28",x"06",x"75",x"D0",x"FA",x"CC",x"98",x"E9",x"76",x"65",x"F9",x"30",x"F7",x"3F",x"10",x"07",x"DE",x"EF",x"1E",x"E9",x"88",x"90",x"E7",x"17",x"84",x"F5",x"DB",x"F4",x"D4",x"51",x"2A",x"60",x"13",x"8A",x"DA",x"2E",x"A7",x"6B",x"4B",x"98",x"A4",x"1C",x"68",x"27",x"43",x"A0",x"76",x"46",x"74",x"B4",x"A6",x"42",x"84",x"4D",x"02",x"29",x"7A",x"5B",x"E9",x"9A",x"A5",x"53",x"57",x"60",x"4C",x"DC",x"68",x"5E",x"D1",x"A4",x"A6",x"D6",x"86",x"0A",x"84",x"E9",x"2C",x"CD",x"4C",x"E6",x"68",x"5E",x"10",x"37",x"28",x"98",x"A0",x"08",x"7F",x"F7",x"F0",x"1D",x"EE",x"4C",x"45",x"82",x"E6",x"0B",x"B3",x"65",x"43",x"85",x"8A",x"AB",x"11",x"68",x"EB",x"22",x"88",x"46",x"D9",x"90",x"03",x"DA",x"44",x"6A",x"66",x"2E",x"88",x"65",x"F4",x"C6",x"10",x"6C",x"37",x"47",x"30",x"02",x"4B",x"18",x"8E",x"0A",x"22",x"78",x"65",x"0B",x"94",x"AB",x"46",x"E8",x"0C",x"C8",x"0B",x"E3",x"8A",x"11",x"DD",x"73",x"35",x"4C",x"FF",x"DE",x"61",x"A2",x"5A",x"DD",x"ED",x"76",x"7F",x"99",x"07",x"19",x"77",x"F7",x"A9",x"12",x"2F",x"BD",x"EE",x"C8",x"76",x"DB",x"60",x"6C",x"0C",x"0D",x"36",x"A9",x"94",x"01",x"4C",x"7B",x"69",x"9F",x"99",x"9E",x"A4",x"9D",x"54",x"3C",x"16",x"D2",x"90",x"91",x"C6",x"6C",x"54",x"1A",x"33",x"65",x"D0",x"48",x"D6",x"C4",x"80",x"D8",x"3D",x"D0",x"88",x"5C",x"11",x"69",x"A5",x"5B",x"A9",x"E9",x"28",x"AA",x"31",x"AA",x"58",x"F2",x"C4",x"3D",x"E2",x"3D",x"60",x"92",x"40",x"0C",x"FE",x"93",x"85",x"AC",x"E4",x"44",x"0E",x"84",x"0F",x"B7",x"A1",x"E0",x"01",x"0C",x"EC",x"C9",x"96",x"DE",x"13",x"56",x"31",x"0D",x"03",x"20",x"85",x"E0",x"68",x"2D",x"0A",x"44",x"0E",x"52",x"0E",x"43",x"41",x"C3",x"00",x"21",x"86",x"9B",x"A2",x"4E",x"46",x"05",x"47",x"04",x"66",x"97",x"6A",x"E2",x"2A",x"A6",x"39",x"69",x"78",x"AF",x"C1",x"10",x"D4",x"18",x"BC",x"84",x"12",x"48",x"ED",x"06",x"1E",x"41",x"0B",x"88",x"AE",x"EF",x"0A",x"A4",x"12",x"77",x"74",x"37",x"88",x"68",x"6C",x"B3",x"4C",x"47",x"64",x"DD",x"8A",x"43",x"48",x"8A",x"7D",x"04",x"8A",x"C1",x"CC",x"15",x"45",x"E4",x"86",x"13",x"84",x"4E",x"5D",x"A4",x"93",x"14",x"47",x"53",x"13",x"98",x"05",x"AA",x"92",x"04",x"34",x"3E",x"99",x"75",x"54",x"1C",x"E7",x"1C",x"E1",x"23",x"14",x"A8",x"D4",x"6E",x"5B",x"35",x"07",x"25",x"34",x"82",x"CD",x"84",x"56",x"D9",x"91",x"0C",x"E6",x"09",x"7A",x"F7",x"45",x"11",x"2D",x"14",x"6B",x"12",x"B6",x"20",x"3F",x"64",x"A8",x"9F",x"72",x"27",x"94",x"68",x"97",x"4C",x"C5",x"12",x"F0",x"A7",x"F5",x"2E",x"31",x"F1",x"A5",x"12",x"D0",x"04",x"F9",x"9D",x"98",x"B5",x"0C",x"24",x"AA",x"61",x"88",x"FC",x"24",x"CF",x"D1",x"46",x"0C",x"AA",x"D5",x"F0",x"10",x"F4",x"DF",x"C0",x"A9",x"A6",x"DB",x"B0",x"03",x"5D",x"FF",x"25",x"01",x"60",x"D6",x"29",x"23",x"EA",x"4E",x"0C",x"F0",x"08",x"E4",x"64",x"F9",x"F6",x"C7",x"E8",x"D0",x"F4",x"98",x"60",x"FB",x"25",x"85",x"9C",x"0C",x"86",x"0D",x"FF",x"E3",x"B0",x"14",x"20",x"D8",x"62",x"5E",x"8D",x"06",x"24",x"81",x"69",x"80",x"B7",x"2E",x"EC",x"E6",x"E7",x"CD",x"E8",x"A5",x"0C",x"EE",x"A6",x"0D",x"60",x"4F",x"38",x"B3",x"88",x"48",x"C8",x"8A",x"E2",x"19",x"71",x"1B",x"AD",x"AA",x"AC",x"DA",x"98",x"49",x"FF",x"38",x"65",x"7E",x"85",x"0D",x"B0",x"75",x"C6",x"03",x"DD",x"42",x"E0",x"65",x"E8",x"26",x"E5",x"27",x"00",x"24",x"60",x"7B",x"FB",x"BB",x"62",x"CB",x"1B",x"D4",x"2E",x"B3",x"03",x"DA",x"EA",x"10",x"E0",x"A0",x"01",x"DE",x"D5",x"01",x"D0",x"BA",x"DE",x"A2",x"83",x"10",x"86",x"11",x"F6",x"50",x"AA",x"D3",x"B8",x"6B",x"6F",x"CE",x"0B",x"60",x"B5",x"A1",x"3B",x"A0",x"10",x"A6",x"ED",x"11",x"F0",x"1F",x"77",x"41",x"26",x"24",x"AA",x"6D",x"A5",x"D9",x"8A",x"11",x"90",x"08",x"85",x"F5",x"05",x"2B",x"93",x"AA",x"2D",x"8A",x"D9",x"E4",x"4B",x"22",x"06",x"0A",x"26",x"0B",x"2A",x"B0",x"7F",x"C5",x"1D",x"90",x"75",x"E5",x"10",x"3D",x"E9",x"88",x"D0",x"EE",x"85",x"04",x"60",x"FE",x"05",x"7A",x"90",x"5E",x"4A",x"A0",x"07",x"ED",x"95",x"69",x"BA",x"71",x"32",x"0D",x"2E",x"8F",x"63",x"CB",x"B0",x"86",x"DA",x"05",x"0B",x"68",x"07",x"A9",x"D6",x"FF",x"15",x"D0",x"0D",x"A5",x"0A",x"F2",x"18",x"21",x"61",x"0F",x"8A",x"6D",x"59",x"5A",x"4C",x"98",x"64",x"48",x"D0",x"C6",x"C4",x"35",x"96",x"CB",x"A0",x"46",x"71",x"E5",x"6D",x"CD",x"C8",x"B1",x"6C",x"8D",x"72",x"D6",x"91",x"CD",x"91",x"02",x"5D",x"EA",x"17",x"5F",x"AD",x"6D",x"5E",x"AE",x"6E",x"79",x"60",x"20",x"FA",x"AF",x"B0",x"A5",x"4A",x"69",x"03",x"AA",x"BD",x"5A",x"3F",x"B5",x"02",x"F0",x"40",x"F7",x"C9",x"FF",x"90",x"E9",x"20",x"4C",x"14",x"5E",x"A0",x"00",x"B1",x"FF",x"A8",x"0A",x"8A",x"86",x"B8",x"D2",x"3A",x"48",x"20",x"B7",x"FF",x"4A",x"7D",x"1E",x"68",x"D6",x"B0",x"A3",x"0E",x"5A",x"02",x"1A",x"0F",x"5A",x"0C",x"DF",x"A7",x"E6",x"0D",x"D0",x"DB",x"20",x"CC",x"FF",x"7F",x"D6",x"8D",x"89",x"7F",x"A5",x"0E",x"A6",x"0F",x"FE",x"60",x"68",x"04",x"57",x"C2",x"10",x"4C",x"4C",x"5E",x"5A",x"91",x"0A",x"EB",x"79",x"85",x"0B",x"A9",x"F4",x"00",x"A8",x"A2",x"06",x"F0",x"3F",x"6A",x"FB",x"E6",x"CC",x"0B",x"CA",x"BB",x"F6",x"C0",x"29",x"F0",x"05",x"91",x"0A",x"FE",x"C8",x"D0",x"F7",x"60",x"50",x"F8",x"5F",x"15",x"65",x"47",x"95",x"90",x"C6",x"72",x"C1",x"06",x"21",x"34",x"6D",x"13",x"B3",x"23",x"31",x"A2",x"0E",x"E5",x"CB",x"B6",x"D1",x"D1",x"F0",x"23",x"2F",x"61",x"F6",x"AB",x"EF",x"C4",x"BC",x"15",x"EF",x"DC",x"75",x"6A",x"27",x"1E",x"2C",x"EB",x"4C",x"2F",x"41",x"17",x"2C",x"92",x"B9",x"8C",x"D0",x"D4",x"9B",x"64",x"51",x"59",x"7E",x"87",x"1A",x"F4",x"92",x"45",x"84",x"58",x"FB",x"A2",x"4C",x"6C",x"73",x"53",x"6C",x"1B",x"6D",x"00",x"25",x"2E",x"40",x"25",x"0B",x"5E",x"11",x"B7",x"B0",x"66",x"42",x"62",x"7A",x"6E",x"6B",x"DD",x"6F",x"A4",x"67",x"72",x"8B",x"6D",x"36",x"0D",x"2A",x"23",x"70",x"17",x"B9",x"F0",x"DE",x"EC",x"49",x"2D",x"8B",x"CB",x"16",x"A2",x"24",x"EC",x"6D",x"77",x"5E",x"97",x"40",x"D1",x"64",x"57",x"5B",x"28",x"3F",x"30",x"43",x"8C",x"49",x"A0",x"EB",x"54",x"01",x"41",x"42",x"93",x"BC",x"CB",x"0C",x"D7",x"09",x"73",x"62",x"61",x"A6",x"6B",x"75",x"9E",x"64",x"C4",x"C5",x"29",x"D4",x"80",x"E3",x"69",x"DA",x"30",x"C9",x"04",x"11",x"F2",x"CF",x"61",x"8F",x"67",x"33",x"DA",x"EE",x"61",x"89",x"63",x"D1",x"61",x"0B",x"2E",x"76",x"92",x"52",x"63",x"F7",x"DC",x"C8",x"72",x"63",x"F4",x"AA",x"50",x"02",x"21",x"A5",x"95",x"22",x"0C",x"16",x"6C",x"E9",x"4A",x"F2",x"79",x"38",x"46",x"57",x"64",x"06",x"5B",x"CF",x"DE",x"C4",x"EC",x"54",x"73",x"11",x"9D",x"28",x"26",x"D0",x"01",x"4A",x"0C",x"68",x"B4",x"48",x"CB",x"D8",x"44",x"1F",x"C0",x"9A",x"2B",x"F4",x"51",x"54",x"35",x"A1",x"22",x"2F",x"8A",x"98",x"9C",x"0F",x"95",x"21",x"B2",x"45",x"DE",x"E4",x"49",x"64",x"26",x"67",x"4E",x"4E",x"65",x"5A",x"4C",x"78",x"25",x"68",x"88",x"AD",x"32",x"66",x"FA",x"E6",x"01",x"4E",x"B2",x"F4",x"BA",x"50",x"52",x"87",x"8C",x"5D",x"76",x"1D",x"26",x"2D",x"70",x"ED",x"81",x"2D",x"87",x"15",x"2C",x"32",x"C4",x"64",x"73",x"5D",x"8F",x"B9",x"B3",x"09",x"D4",x"D7",x"12",x"A8",x"8A",x"73",x"60",x"12",x"41",x"38",x"67",x"A7",x"40",x"65",x"56",x"9B",x"3D",x"12",x"D4",x"43",x"A4",x"22",x"2C",x"99",x"4B",x"B0",x"CD",x"93",x"A4",x"09",x"6D",x"15",x"2E",x"62",x"EE",x"80",x"73",x"12",x"4C",x"DE",x"EB",x"73",x"FB",x"4B",x"B3",x"65",x"4B",x"45",x"D8",x"59",x"6F",x"39",x"30",x"5A",x"8C",x"BA",x"E4",x"26",x"D8",x"E4",x"76",x"99",x"DD",x"3F",x"6D",x"09",x"11",x"8D",x"64",x"62",x"75",x"A3",x"1A",x"25",x"D5",x"4D",x"B3",x"0B",x"60",x"71",x"6D",x"CF",x"D4",x"53",x"79",x"73",x"F8",x"CA",x"6D",x"56",x"A3",x"44",x"80",x"18",x"4A",x"80",x"D2",x"30",x"73",x"29",x"2D",x"D8",x"C1",x"5C",x"74",x"6B",x"A6",x"03",x"35",x"C5",x"68",x"AD",x"33",x"29",x"B2",x"CB",x"33",x"E3",x"00",x"13",x"37",x"69",x"A5",x"64",x"52",x"36",x"24",x"6E",x"87",x"28",x"94",x"63",x"94",x"68",x"2E",x"8F",x"54",x"8A",x"7A",x"B4",x"7B",x"CE",x"E7",x"7A",x"B6",x"AC",x"56",x"F3",x"48",x"2B",x"44",x"46",x"8E",x"50",x"AB",x"A1",x"41",x"8E",x"6C",x"58",x"A1",x"B4",x"0A",x"5D",x"E4",x"C7",x"62",x"B5",x"25",x"0E",x"7A",x"85",x"EC",x"08",x"62",x"3A",x"E8",x"00",x"4F",x"A0",x"76",x"D6",x"64",x"69",x"39",x"28",x"31",x"8F",x"95",x"45",x"78",x"EE",x"E2",x"18",x"6D",x"CB",x"D6",x"E7",x"01",x"57",x"28",x"65",x"81",x"4A",x"61",x"F6",x"C6",x"15",x"74",x"8A",x"20",x"8F",x"27",x"73",x"53",x"D1",x"71",x"3A",x"CE",x"79",x"70",x"1E",x"65",x"4D",x"8D",x"78",x"CE",x"11",x"A4",x"65",x"8A",x"55",x"3A",x"7C",x"55",x"D6",x"35",x"CA",x"23",x"E5",x"6D",x"A4",x"62",x"85",x"45",x"E7",x"09",x"DB",x"5A",x"88",x"E8",x"4E",x"09",x"30",x"E1",x"28",x"49",x"10",x"6B",x"35",x"44",x"73",x"6C",x"E6",x"45",x"29",x"5B",x"41",x"6B",x"52",x"02",x"70",x"3D",x"9A",x"D1",x"8A",x"15",x"7A",x"3C",x"06",x"2E",x"C0",x"ED",x"22",x"68",x"7C",x"5B",x"CA",x"41",x"A5",x"CE",x"B9",x"4B",x"27",x"71",x"8A",x"2E",x"4C",x"76",x"E2",x"E8",x"42",x"D4",x"62",x"53",x"E6",x"31",x"02",x"99",x"45",x"D9",x"73",x"B1",x"AE",x"46",x"89",x"D2",x"59",x"67",x"BB",x"72",x"15",x"31",x"42",x"7A",x"5A",x"49",x"61",x"94",x"C0",x"4E",x"B7",x"1A",x"54",x"94",x"1D",x"56",x"24",x"B9",x"56",x"C8",x"4A",x"90",x"62",x"75",x"73",x"FC",x"95",x"5C",x"57",x"1B",x"1C",x"52",x"E3",x"7C",x"44",x"66",x"DB",x"5E",x"16",x"79",x"11",x"D8",x"60",x"43",x"75",x"37",x"E4",x"36",x"5B",x"F7",x"70",x"14",x"8E",x"D2",x"4B",x"6E",x"2A",x"A9",x"5C",x"5B",x"3A",x"2B",x"D3",x"47",x"35",x"76",x"A5",x"EF",x"FE",x"4E",x"10",x"46",x"98",x"72",x"7A",x"A1",x"36",x"37",x"64",x"69",x"4F",x"BD",x"04",x"7B",x"28",x"84",x"23",x"29",x"1B",x"D3",x"2D",x"11",x"20",x"46",x"D5",x"44",x"73",x"00",x"06",x"21",x"45",x"E7",x"39",x"25",x"88",x"4D",x"CE",x"D1",x"EA",x"AA",x"44",x"29",x"8B",x"B3",x"57",x"71",x"33",x"55",x"03",x"40",x"3D",x"2C",x"6F",x"4A",x"F3",x"72",x"B6",x"6F",x"6F",x"70",x"D1",x"75",x"9D",x"61",x"9E",x"67",x"90",x"2F",x"4A",x"94",x"5C",x"9A",x"62",x"85",x"A6",x"48",x"AA",x"20",x"A4",x"63",x"6F",x"97",x"9C",x"C8",x"75",x"65",x"87",x"ED",x"4B",x"4C",x"B4",x"51",x"2B",x"62",x"D5",x"56",x"96",x"78",x"59",x"54",x"48",x"71",x"FF",x"47",x"00",x"1B",x"96",x"78",x"FC",x"B1",x"2D",x"77",x"B3",x"56",x"89",x"6E",x"00",x"DB",x"6D",x"65",x"67",x"61",x"AF",x"64",x"90",x"38",x"93",x"FD",x"66",x"A8",x"2E",x"78",x"61",x"4D",x"6B",x"9D",x"00",x"42",x"E1",x"DE",x"43",x"48",x"6E",x"D5",x"4F",x"44",x"45",x"EE",x"69",x"74",x"42",x"18",x"78",x"74",x"D2",x"C6",x"6E",x"61",x"DE",x"6C",x"CB",x"49",x"58",x"66",x"EC",x"42",x"52",x"46",x"A5",x"54",x"6D",x"61",x"74",x"17",x"72",x"29",x"1B",x"B4",x"73",x"49",x"A5",x"31",x"0A",x"30",x"2F",x"00",x"BB",x"CA",x"2A",x"E2",x"47",x"53",x"4A",x"7A",x"74",x"B6",x"2D",x"0B",x"88",x"5C",x"95",x"5D",x"7F",x"3D",x"2D",x"24",x"40",x"2F",x"04",x"25",x"90",x"D2",x"3B",x"0F",x"09",x"00",x"02",x"7C",x"00",x"C0",x"EB",x"12",x"2D",x"60",x"58",x"77",x"B0",x"32",x"34",x"73",x"E4",x"A9",x"28",x"15",x"29",x"C2",x"5D",x"50",x"59",x"B9",x"D1",x"47",x"48",x"9D",x"DA",x"89",x"31",x"37",x"BD",x"65",x"30",x"0B",x"32",x"5A",x"50",x"49",x"55",x"5D",x"47",x"16",x"3F",x"79",x"A5",x"2D",x"42",x"AC",x"4F",x"50",x"48",x"5A",x"4E",x"D4",x"B3",x"43",x"A7",x"64",x"00",x"36",x"92",x"02",x"AA",x"15",x"C7",x"6F",x"6D",x"31",x"48",x"41",x"53",x"E2",x"DD",x"07",x"43",x"55",x"5D",x"45",x"44",x"C3",x"B6",x"56",x"6F",x"52",x"1F",x"49",x"3F",x"C0",x"02",x"20",x"00",x"30",x"F0",x"49",x"92",x"CB",x"6E",x"4F",x"59",x"EE",x"25",x"B3",x"73",x"E5",x"7D",x"46",x"6F",x"75",x"6E",x"EF",x"72",x"66",x"69",x"D7",x"3A",x"BA",x"20",x"01",x"46",x"2E",x"28",x"60",x"3F",x"EF",x"48",x"6E",x"FD",x"0F",x"E0",x"80",x"81",x"6B",x"DA",x"D6",x"DB",x"B4",x"50",x"92",x"14",x"EB",x"D2",x"55",x"2E",x"4E",x"3B",x"AB",x"D1",x"3D",x"76",x"35",x"EC",x"DD",x"0A",x"35",x"2B",x"45",x"52",x"4D",x"DD",x"E4",x"20",x"55",x"DE",x"53",x"4C",x"68",x"9E",x"59",x"00",x"F7",x"B6",x"A9",x"24",x"31",x"51",x"53",x"66",x"70",x"65",x"A1",x"64",x"43",x"3D",x"01",x"20",x"4B",x"C5",x"42",x"2F",x"93",x"00",x"56",x"C8",x"15",x"DF",x"9C",x"79",x"32",x"31",x"66",x"92",x"C1",x"1C",x"44",x"08",x"4D",x"5D",x"78",x"69",x"47",x"75",x"6D",x"3B",x"72",x"AD",x"64",x"A2",x"61",x"62",x"6C",x"0F",x"AD",x"65",x"63",x"74",x"75",x"10",x"61",x"73",x"DA",x"3A",x"57",x"D9",x"69",x"74",x"EA",x"A8",x"65",x"14",x"8A",x"6F",x"72",x"8E",x"40",x"20",x"06",x"38",x"24",x"47",x"56",x"91",x"02",x"4D",x"69",x"42",x"17",x"53",x"15",x"43",x"B6",x"52",x"72",x"7B",x"46",x"4F",x"55",x"B7",x"F6",x"2E",x"00",x"30",x"31",x"32",x"33",x"FE",x"3C",x"36",x"37",x"38",x"EF",x"39",x"C1",x"C2",x"C3",x"C4",x"C5",x"C6",x"2D",x"FF",x"32",x"31",x"87",x"37",x"0E",x"33",x"36",x"34",x"38",x"BB",x"7B",x"0C",x"9D",x"09",x"0A",x"10",x"40",x"50",x"A0",x"D0",x"FF",x"27",x"A6",x"93",x"7A",x"2A",x"00",x"30",x"33",x"41",x"40",x"48",x"44",x"14",x"68",x"C0",x"11",x"01",x"F1",x"53",x"01",x"C0",x"1C",x"06",x"22",x"68",x"05",x"16",x"86",x"66",x"09",x"9D",x"C5",x"80",x"C8",x"55",x"25",x"1B",x"E0",x"22",x"68",x"4E",x"03",x"64",x"E6",x"03",x"B6",x"95",x"01",x"05",x"74",x"CB",x"05",x"2C",x"08",x"07",x"09",x"04",x"14",x"FA",x"15",x"06",x"D1",x"16",x"17",x"6B",x"18",x"0D",x"19",x"9D",x"1A",x"03",x"1B",x"1E",x"1C",x"0B",x"1D",x"06",x"1E",x"FD",x"1F",x"0D",x"20",x"E9",x"21",x"35",x"22",x"07",x"27",x"01",x"31",x"FA",x"03",x"32",x"0E",x"33",x"1F",x"34",x"08",x"3C",x"06",x"3D",x"FD",x"3E",x"01",x"3F",x"EA",x"09",x"40",x"4F",x"41",x"0E",x"42",x"07",x"43",x"7F",x"46",x"06",x"47",x"7A",x"48",x"08",x"49",x"EB",x"03",x"4A",x"04",x"4B",x"3F",x"07",x"4E",x"0B",x"EC",x"2A",x"42",x"49",x"C5",x"53",x"54",x"D1",x"27",x"4D",x"94",x"30",x"87",x"FF",x"85",x"26",x"39",x"EB",x"58",x"90",x"9F",x"56",x"72",x"31",x"FC",x"08",x"B2",x"E2",x"DD",x"CA",x"78",x"C6",x"62",x"E8",x"0F",x"B8",x"F8",x"20",x"2A",x"02",x"A3",x"1B",x"11",x"06",x"01",x"07",x"28",x"29",x"6D",x"CA",x"66",x"62",x"61",x"97",x"E1",x"21",x"4B",x"46",x"41",x"54",x"33",x"32",x"3E",x"20",x"B0",x"0E",x"1F",x"BE",x"77",x"7C",x"AC",x"22",x"C0",x"FF",x"74",x"0B",x"56",x"B4",x"0E",x"BB",x"07",x"00",x"FF",x"10",x"AC",x"5E",x"5B",x"F0",x"32",x"E4",x"8F",x"16",x"CD",x"19",x"EB",x"FE",x"7E",x"03",x"8B",x"48",x"59",x"D7",x"50",x"A0",x"42",x"A1",x"4F",x"A0",x"8A",x"56",x"16",x"30",x"2E",x"1A",x"31",x"74",x"6F",x"0D",x"3F",x"4E",x"4F",x"7F",x"47",x"90",x"53",x"34",x"CF",x"87",x"24",x"5B",x"63",x"65",x"E6",x"5D",x"59",x"32",x"2C",x"36",x"D7",x"C3",x"38",x"38",x"35",x"31",x"E4",x"30",x"9F",x"50",x"6E",x"43",x"2C",x"0B",x"53",x"94",x"0C",x"20",x"34",x"B3",x"4F",x"50",x"16",x"DD",x"36",x"63",x"99",x"54",x"2C",x"44",x"E9",x"53",x"4B",x"B4",x"B4",x"1A",x"D5",x"42",x"4C",x"BA",x"43",x"4F",x"4D",x"50",x"55",x"7E",x"45",x"53",x"56",x"4E",x"44",x"D9",x"54",x"52",x"D3",x"59",x"20",x"47",x"24",x"49",x"4E",x"77",x"0B",x"6A",x"52",x"45",x"41",x"44",x"59",x"2E",x"FD",x"0D",x"0A",x"00",x"3F",x"0C",x"34",x"20",x"F8",x"53",x"0F",x"BB",x"08",x"0F",x"45",x"61",x"53",x"AE",x"93",x"4A",x"BE",x"30",x"38",x"02",x"03",x"0E",x"10",x"4D",x"91",x"D1",x"2B",x"72",x"45",x"4D",x"2E",x"C9",x"21",x"4D",x"45",x"47",x"41",x"36",x"35",x"FE",x"59",x"53",x"D1",x"30",x"A0",x"80",x"A1",x"08",x"9C",x"B2",x"4B",x"46",x"ED",x"74",x"CF",x"2A",x"06",x"32",x"32",x"3E",x"32",x"90",x"D1",x"1A",x"E2",x"6A",x"6E",x"8A",x"33",x"06",x"47",x"9B",x"34",x"1B",x"4D",x"B3",x"69",x"B4",x"05",x"51",x"89",x"EC",x"46",x"26",x"B2",x"09",x"63",x"85",x"04",x"4A",x"54",x"00",x"65",x"09",x"D5",x"D3",x"58",x"52",x"04",x"03",x"02",x"07",x"F5",x"06",x"08",x"7F",x"75",x"CF",x"28",x"C6",x"20",x"61",x"02",x"01",x"D7",x"72",x"13",x"B0",x"16",x"86",x"19",x"DE",x"5C",x"4F",x"51",x"46",x"87",x"47",x"95",x"9E",x"4D",x"4A",x"8E",x"4E",x"2F",x"57",x"B2",x"88",x"B9",x"C6",x"8D",x"56",x"6C",x"8C",x"59",x"79",x"E9",x"20",x"A1",x"E8",x"E6",x"D0",x"E8",x"60",x"01",x"1E",x"02",x"F4",x"50",x"80",x"03",x"22",x"11",x"8C",x"6C",x"01",x"0A",x"00",x"A0",x"02",x"F0",x"F0",x"07",x"A9",x"C8",x"AF",x"4C",x"A4",x"38",x"5B",x"60",x"A2",x"19",x"B5",x"02",x"9D",x"77",x"79",x"FF",x"CA",x"10",x"F8",x"6F",x"00",x"A2",x"D0",x"85",x"02",x"86",x"FD",x"03",x"9B",x"0E",x"D2",x"56",x"90",x"91",x"15",x"04",x"D6",x"BE",x"79",x"A9",x"05",x"F5",x"A2",x"03",x"A0",x"97",x"20",x"BA",x"96",x"4C",x"C0",x"FF",x"B7",x"79",x"3E",x"89",x"C8",x"84",x"BB",x"B3",x"22",x"A2",x"99",x"89",x"50",x"67",x"4D",x"84",x"3B",x"AB",x"22",x"A2",x"19",x"A1",x"10",x"AB",x"91",x"19",x"11",x"91",x"B9",x"87",x"3A",x"99",x"E6",x"07",x"88",x"D0",x"F7",x"18",x"AA",x"98",x"29",x"0F",x"99",x"68",x"03",x"F0",x"0C",x"8A",x"79",x"67",x"03",x"99",x"68",x"03",x"A5",x"9F",x"79",x"9B",x"03",x"99",x"9C",x"03",x"A9",x"01",x"85",x"9F",x"A9",x"78",x"20",x"00",x"01",x"4A",x"AA",x"F0",x"09",x"08",x"06",x"9F",x"38",x"6A",x"CA",x"D0",x"F9",x"28",x"6A",x"99",x"34",x"03",x"30",x"05",x"A5",x"9F",x"86",x"9F",x"24",x"8A",x"C8",x"C0",x"34",x"D0",x"C1",x"A0",x"C9",x"8A",x"4C",x"9C",x"01",x"22",x"00",x"79",x"69",x"80",x"0A",x"10",x"0F",x"06",x"FD",x"D0",x"08",x"48",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"68",x"2A",x"30",x"F1",x"70",x"01",x"60",x"38",x"85",x"A7",x"AD",x"29",x"01",x"D0",x"06",x"CE",x"2A",x"01",x"8E",x"E7",x"DB",x"CE",x"29",x"01",x"AD",x"91",x"39",x"60",x"20",x"1A",x"01",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"66",x"A8",x"CA",x"06",x"FD",x"D0",x"06",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"E8",x"90",x"F3",x"F0",x"E1",x"E0",x"11",x"B0",x"51",x"BD",x"33",x"03",x"20",x"00",x"01",x"7D",x"67",x"03",x"85",x"9E",x"AA",x"24",x"A8",x"10",x"09",x"70",x"07",x"A9",x"00",x"20",x"05",x"01",x"D0",x"25",x"A9",x"F1",x"E0",x"03",x"B0",x"03",x"BD",x"A2",x"01",x"B8",x"20",x"05",x"01",x"18",x"AA",x"BD",x"34",x"03",x"20",x"00",x"01",x"7D",x"68",x"03",x"85",x"AE",x"A5",x"A7",x"7D",x"9C",x"03",x"65",x"FF",x"85",x"AF",x"A6",x"9E",x"B1",x"AE",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"CA",x"D0",x"F1",x"86",x"A7",x"F0",x"99",x"4C",x"0D",x"08",x"CC",x"F2",x"01",x"00",x"0B",x"9C",x"F0",x"03",x"9E",x"32",x"30",x"36",x"31",x"7E",x"60",x"10",x"7F",x"4E",x"8D",x"D5",x"29",x"F8",x"09",x"06",x"F6",x"85",x"01",x"BA",x"8E",x"CF",x"9A",x"9D",x"E8",x"82",x"C6",x"6C",x"77",x"B1",x"1D",x"48",x"C8",x"AD",x"28",x"7F",x"19",x"BD",x"77",x"79",x"5F",x"02",x"BD",x"FB",x"68",x"97",x"85",x"50",x"52",x"4F",x"50",x"2E",x"4D",x"36",x"35",x"55",x"2E",x"4E",x"41",x"4D",x"45",x"3D",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"46",x"44",x"49",x"53",x"4B",x"2B",x"46",x"4F",x"52",x"4D",x"41",x"54",x"20",x"55",x"54",x"49",x"4C",x"49",x"54",x"59",x"4D",x"36",x"35",x"55",x"4B",x"45",x"59",x"42",x"4F",x"41",x"52",x"44",x"20",x"54",x"45",x"53",x"54",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"95",x"01",x"0D",x"08",x"44",x"56",x"05",x"58",x"01",x"08",x"0B",x"08",x"37",x"01",x"9E",x"32",x"30",x"36",x"31",x"00",x"00",x"00",x"BA",x"BD",x"9A",x"08",x"9D",x"FC",x"00",x"CA",x"D0",x"F7",x"A0",x"35",x"4C",x"4C",x"08",x"DD",x"55",x"2E",x"4E",x"7F",x"4D",x"3D",x"AD",x"4B",x"59",x"BF",x"42",x"4F",x"41",x"52",x"44",x"20",x"7F",x"45",x"53",x"54",x"00",x"3D",x"09",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B9",x"42",x"09",x"99",x"E6",x"07",x"88",x"D0",x"F7",x"18",x"AA",x"98",x"29",x"0F",x"99",x"68",x"03",x"F0",x"0C",x"8A",x"79",x"67",x"03",x"99",x"68",x"03",x"A5",x"9F",x"79",x"9B",x"03",x"99",x"9C",x"03",x"A9",x"01",x"85",x"9F",x"A9",x"78",x"20",x"00",x"01",x"4A",x"AA",x"F0",x"09",x"08",x"06",x"9F",x"38",x"6A",x"CA",x"D0",x"F9",x"28",x"6A",x"99",x"34",x"03",x"30",x"05",x"A5",x"9F",x"86",x"9F",x"24",x"8A",x"C8",x"C0",x"34",x"D0",x"C1",x"A0",x"54",x"8A",x"4C",x"9C",x"01",x"02",x"00",x"08",x"69",x"80",x"0A",x"10",x"0F",x"06",x"FD",x"D0",x"08",x"48",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"68",x"2A",x"30",x"F1",x"70",x"01",x"60",x"38",x"85",x"A7",x"AD",x"29",x"01",x"D0",x"06",x"CE",x"2A",x"01",x"8E",x"E7",x"DB",x"CE",x"29",x"01",x"AD",x"4C",x"08",x"60",x"20",x"1A",x"01",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"66",x"A8",x"CA",x"06",x"FD",x"D0",x"06",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"E8",x"90",x"F3",x"F0",x"E1",x"E0",x"11",x"B0",x"51",x"BD",x"33",x"03",x"20",x"00",x"01",x"7D",x"67",x"03",x"85",x"9E",x"AA",x"24",x"A8",x"10",x"09",x"70",x"07",x"A9",x"00",x"20",x"05",x"01",x"D0",x"25",x"A9",x"F1",x"E0",x"03",x"B0",x"03",x"BD",x"A2",x"01",x"B8",x"20",x"05",x"01",x"18",x"AA",x"BD",x"34",x"03",x"20",x"00",x"01",x"7D",x"68",x"03",x"85",x"AE",x"A5",x"A7",x"7D",x"9C",x"03",x"65",x"FF",x"85",x"AF",x"A6",x"9E",x"B1",x"AE",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"CA",x"D0",x"F1",x"86",x"A7",x"F0",x"99",x"4C",x"0E",x"08",x"CC",x"F2",x"01",x"00",x"0B",x"08",x"0A",x"DC",x"9E",x"B5",x"30",x"36",x"32",x"0E",x"00",x"78",x"F1",x"47",x"92",x"53",x"70",x"2F",x"3D",x"41",x"85",x"A9",x"A7",x"00",x"11",x"77",x"20",x"D6",x"21",x"80",x"CE",x"6F",x"D0",x"A9",x"FF",x"F6",x"15",x"5B",x"8D",x"16",x"D6",x"4C",x"FF",x"08",x"5A",x"52",x"4F",x"50",x"6F",x"36",x"35",x"50",x"52",x"4F",x"50",x"2E",x"4D",x"36",x"35",x"55",x"2E",x"4E",x"41",x"4D",x"45",x"3D",x"4B",x"45",x"59",x"42",x"4F",x"41",x"52",x"44",x"20",x"54",x"45",x"53",x"54",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");

begin  -- behavioural

  process(clka)
  begin

    --report "COLOURRAM: A Reading from $" & to_hstring(unsigned(addra))
    --  & " = $" & to_hstring(ram(to_integer(unsigned(addra))));
    if(rising_edge(Clka)) then 
      if ena='1' then
        if(wea="1") then
          ram(to_integer(unsigned(addra(14 downto 0)))) := dina;
          report "COLOURRAM: A writing to $" & to_hstring(unsigned(addra))
            & " = $" & to_hstring(dina);
            douta <= dina;
          else
            douta <= ram(to_integer(unsigned(addra(14 downto 0))));            
        end if;
      end if;
    end if;
  end process;

  process (clkb)
  begin
    if(rising_edge(Clkb)) then 
      if(web="1") then
--        ram(to_integer(unsigned(addrb))) <= dinb;
      end if;
      doutb <= ram(to_integer(unsigned(addrb(14 downto 0))));
    end if;
  end process;

end behavioural;
