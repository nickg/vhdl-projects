-- *********************************************************************/ 
-- Copyright 2006 Actel Corporation.  All rights reserved.
-- IP Solutions Group
--  
-- File:  EDAC NETLIST
--     
-- Description: EDAC
--                
--
-- Rev: 1.0  01Jul02 HC  : Initial Code  
-- Rev: 1.3  17May06 IPB : Fixed Simultanous read/write SARS
-- Rev: 1.4  01Jun06 IPB : Removed W2R port
-- Rev: 1.5  06Jun06 IPB : fixed SLOWDOWN issue SAR	56406
--
-- Notes:
--
--
-- *********************************************************************/ 
--
--
--
library IEEE,axcelerator;

use IEEE.std_logic_1164.all;
use axcelerator.components.all;

package CONV_PACK_edaci is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_edaci;

library IEEE,axcelerator;

use IEEE.std_logic_1164.all;
use axcelerator.components.all;

use work.CONV_PACK_edaci.all;

entity edaci is

   port( waddr, raddr : in std_logic_vector (11 downto 0);  wdata : in 
         std_logic_vector (28 downto 0);  rdata : out std_logic_vector (28 
         downto 0);  tmout : in std_logic_vector (41 downto 0);  rds : in 
         std_logic_vector (3 downto 0);  wp : in std_logic_vector (6 downto 0);
         rp : out std_logic_vector (6 downto 0);  caddr, axwaddr, axraddr : out
         std_logic_vector (11 downto 0);  axwdata : out std_logic_vector (35 
         downto 0);  axrdata : in std_logic_vector (35 downto 0);  clk, we, re,
         rstn, stop_scrub, bypass : in std_logic;  slowdown, scrub_corrected, 
         error, scrub_done, tmoutflg, correctable, axwe, axre : out std_logic);

end edaci;

architecture SYN_DEF_ARCH of edaci is

signal VXXXXXXXX, XXXDXXXXXXXXXXXXXXXXXX, XXDDXXXXXQ, XXDXXXXXX, XXDDXXXXXJ, 
   XXYPXXXXXX, XXYPXXXXXXF, XXDDXXXXXL, XXDDXXXXX, XXXXXXDXXXX, XXDDXXXXXW, 
   XXDDXXXXXXF, XXXXXXXXXXXXXXDX, XXXXXXXXXLXXF, XXDDXXXXXX, XXYPXXXXXXH, 
   XXDDXXXXXF, XXDDXXXXXV, XXDDXXXXXK, XXDDXXXXXH, XXDDXXXXXP, XXDXXXXXXXXXX, 
   XXDXXXXXXXXXXF, XXDXXXXXXXXXXH, XXDXXXXXXXXXXXXXX, XXDXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXF, XXDXXXXXXXXXXK, XXDXXXXXXXXXXL, XXDXXXXXXXXXXP, 
   XXDXXXXXXXXXXQ, XXDXXXXXXXXXXV, XXDXXXXXXXXXXW, XXDXXXXXXXX, XXDXXXXXXXXXXFD
   , XXDXXXXXXXXXXFF, XXDXXXXXXXXXXXXXXH, XXDXXXXXXXXXXFH, XXDXXXXXXXXXXFJ, 
   XXDXXXXXXXXXXFK, XXDXXXXXXXXXXFL, XXDXXXXXXXXF, XXDXXXXXXXXXXFP, 
   XXDXXXXXXXXXXFQ, XXDXXXXXXXXXXFV, XXDXXXXXXXXXXFW, XXDXXXXXXXXXXHD, 
   XXDXXXXXXXXXXHF, XXDXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXHH, XXDXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXHJ, XXDXXXXXXXXH, XXDXXXXXXXXXXHK, XXDXXXXXXXXXXHL, 
   XXDXXXXXXXXXXHP, XXDXXXXXXXXXXHQ, XXDXXXXXXXXXXHV, XXDXXXXXXXXXXHW, 
   XXDXXXXXXXXXXJD, XXDXXXXXXXXXXJF, XXDXXXXXXXXXXXXXXL, XXDXXXXXXXXXXJH, 
   XXDXXXXXXXXXXXXXXP, XXDXXXXXXXXXXJJ, XXDXXXXXXXXXXJK, XXDXXXXXXXXXXJL, 
   XXDXXXXXXXXXXJP, XXDXXXXXXXXXXJQ, XXDXXXXXXXXJ, XXDXXXXXXXXXXJV, 
   XXDXXXXXXXXXXJW, XXDXXXXXXXXXXKD, XXDXXXXXXXXXXXDXDXXXXXXXXFV, 
   XXDXXXXXXXXXXXDXDXXXXXXXXFW, XXDXXXXXXXXXXXDXDXXXXXXXXHD, 
   XXDXXXXXXXXXXXDXDXXXXXX, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXDXDXXXXXXF, XXDXXXXXXXXXXXDXDXXXXXXH, 
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXDXDXXXXXXXXHF, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXDXDXXXXXXJ, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXP, XXDXXXXXXXXXXXDXDXXXXXXXXHH, 
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXQ, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXV, 
   XXDXXXXXXXXXXXXXXXDXDX, XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXXXXXXXXDXDX, 
   XXDXXXXXXXXXXXDXDXXXXXXK, XXDXXXXXXXXXXXDXDXXXXXXXXHJ, 
   XXDXXXXXXXXXXXDXDXXXXXXXXHK, XXDXXXXXXXXXXXDXDXXXXXXL, 
   XXDXXXXXXXXXXXDXDXXXXXXP, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXF, XXDXXXXDXXXXXXXXXX, XXDXXXXDXXXXXXXX, 
   XXDXXXXDXXXXXXXXF, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXH, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF
   , XXDXXXXDXXXXXYXXXXXXXXXXXXXJ, XXDXXXXDXXXXXYXXXXXXXXXXXXXK, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXDXXXXXYXXXXXXXXXXXXXL, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXXX, XXDXXXXDXXXXXYXXXXXXXHD, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXP, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH
   , XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF
   , XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, 
   XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXX, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, XXDXXXXDXXXXXYXXXXXXXXXXXXXQ, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXV, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXF, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, XXDXXXXDXXXXXYXXXXXXXXXXXXXW
   , XXDXXXXDXXXXXYXXXXXXXXXXXXXFD, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXFF, XXDXXXXDXXXXXYXXXXXXXXXXXXXFH, 
   XXDXXXXDXXXXXXXXH, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXXXH, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, 
   XXDXXXXDXXXXXYXXXXX, XXDXXXXDXXXXXXXXXXF, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXJ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXK, 
   XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXXXX, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXL, 
   XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXX, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP
   , XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXP, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXFJ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, XXDXXXXDXXXXXYXXXXXF, 
   XXDXXXXDXXXXXYXXXXXH, XXDXXXXDXXXXXXXXJ, XXDXXXXDXXXXXYXXXXXXXXXXXXXFK, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXF, XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ,
   XXDXXXXDXXXXXYXXXXXXXXXXXXXFL, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, XXDXXXXDXXXXXXXXK, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXH,
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, XXDXXXXDXXXXXYXXXXXXXXXXXXXFP, 
   XXDXXXXDXXXXXYXXXXXJ, XXDXXXXDXXXXXYXXXXXK, XXDXXXXDXXXXXYXXXXXXXXXXXXXFQ, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXFV, XXDXXXXDXXXXXYXXXXXXXXXXXXXFW, 
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, XXDXXXXDXXXXXXXXL, 
   XXDXXXXDXXXXXYXXXXXXXXXXXXXHD, XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXDXXXXXXXFLXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, XXDXXXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXX, XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXYXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXXXXXXXXXXXXXXXJW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, XXDXXXXXXXXXXY, XXDXXXXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXXXXXXXKD, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXKF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXJ, XXDXXXXXXXXXXXXXXXXXXXXLXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXFF, XXDXXXXXXXXXXXXXXXXXXXXXXXXKH, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXX, XXDXXXXXXXXXXYXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXFD, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXYXXF, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXP, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXKJ, 
   XXDXXXXXXXXXXXXXXDDXXLXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXQ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXF
   , XXDXXXXXXXXXXXXXXXXXXXXXXQXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXKK, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXJ, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXFF, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXKL, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXX, XXDXXXXXXXXXXXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXKP, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXKQ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXF, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXK, XXDXXXXXXXXXXXXXXXXXXXXXXXXKV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, XXDXXXXXXXXXXXXXXXXXXXXXXXXKW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXFH, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, XXDXXXXXXXXXXXXXXXXXXXXXXXFJ, 
   XXDXXXXXXXXXXXXXXXFH, XXDXXXXXXXXXXXFXXXXLXXDX, XXDXXXXXXXXXXYXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, XXDXXXXXXXXXXXXXXDDXXLXX, 
   XXDXXXXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXXFJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXH, XXDXXXXXXXXXXXXXXXDDXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXQ, 
   XXDXXXXXXXXXXXXXXDDXXXXXFD, XXDXXXXXXXXXXXXXXXXXXXXLXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXL, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXQ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, 
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXV,
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, XXDXXXXXXXXXXXXXXDDXXLXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXV, XXDXXXXXXXXXXYXXJ, XXDXXXXXXXXXXXXXXXFK, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK
   , XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, 
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXLXXXW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFD, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, 
   XXDXXXXXXXXXXXXXXDDXXXXXXXXXX, XXDXXXXXXXXXXXXXXXFL, XXDXXXXXXXXXXXXXXXFP, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFD, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFF, XXDXXXXXXXXXXXXWXX, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXYXXK, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, 
   XXDXXXXXXXXXXXXXXDDXXLXXH, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFD, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFH, 
   XXDXXXXXXXXXXXXXXDDXXLXXJ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFH, XXDXXXXXXXXXXXXXXXXXXXXLXXXFJ, 
   XXDXXXXXXXXXXXXXXXWXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXXXXXLD, 
   XXDXXXXXXXXXXXXXXDDXXXXXFF, XXDXXXXXXXXXXXXXXXWXXXXXXXX, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFH, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFK, 
   XXDXXXXXXXXXXYXXL, XXDXXXXXXXXXXXXXXDDXXLXXX, XXDXXXXXXXXXXXXXXDDXXLXXK, 
   XXDXXXXXXXXXXYXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFK, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFL, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXFP, XXDXXXXXXXXXXXXXXDDXXLXXL, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFJ, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFK, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, XXDXXXXXXXXXXXXXXXXXXXXLXXXFQ, 
   XXDXXXXXXXXXXXXXXDDXXLXXP, XXDXXXXXXXXXXXXXXDDXXXXXFH, XXDXXXXXXXXXXXXXXXFQ,
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXK, XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX, 
   XXDXXXXXXXXXXYXXP, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, XXDXXXXXXXXXXXXXXDDXXXXXFJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXDDXXLXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXL, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXFV, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXFW, 
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXK, XXDXXXXXXXXXXXXXXXFLXX, 
   XXDXXXXXXXXXXXXXXXXXJ, XXDXXXXXXXXXXYXXXH, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFP
   , XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHD, XXDXXXXXXXXXXXXXXXFV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXLF, XXDXXXXXXXXXXXXXXDDXXXXXFK, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXL, XXDXXXXXXXXXXXXXXXFW, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFQ, XXDXXXXXXXXXXXXXXXXXXXXLXXXHH, 
   XXDXXXXXXXXXXXXXXDDXXLXXQ, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFV, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFL, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXP, XXDXXXXXXXXXXXXXXXXXXXXLXXXHJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXDDXXLXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHK, XXDXXXXXXXXXXXXXXDDXXLXXXXXXXF, 
   XXDXXXXXXXXXXXXPXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXHL, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFP, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP, XXDXXXXXXXXXXXXXXXHD, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK,
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXLXXXHP, 
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHQ, XXDXXXXXXXXXXXXXXDDXXLXXW, 
   XXDXXXXXXXXXXXXXXXHF, XXDXXXXXXXXXXXXXXXXXXXXLXXXHV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, XXDXXXXXXXXXXXXXXXHH, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXHW, XXDXXXXXXXXXXYXXQ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFQ, 
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFV, 
   XXDXXXXXXXXXXXXXXDDXXXXXFL, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXQ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXHJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFW, 
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXJD, 
   XXDXXXXXXXXXXXXXXXHK, XXDXXXXXXXXXXXXXXXXXXXXLXXL, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXYXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHD, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHD, XXDXXXXXXXXXXXXXXDDXXLXXXXXXXH, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHF, XXDXXXXXXXXXXXXXXXXXXXXXXXXLH, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, 
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHH, XXDXXXXXXXXXXXXXXXXXXXXXXXXLJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHJ, 
   XXDXXXXXXXXXXXXXDDXXF, XXDXXXXXXXXXXXXXXXHL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXYXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHK, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, XXDXXXXXXXXXXXXXXXXXXXXLXXP, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHH, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXLK, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHL, 
   XXDXXXXXXXXXXXXXXXHP, XXDXXXXXXXXXXXXXXXXXXXXXXXXLL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, 
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, XXDXXXXXXXXXXXXXXXXXXXXXXXXLP, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHJ, XXDXXXXXXXXXXXXXXXXXXXXLXXXJF, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHP, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHK, 
   XXDXXXXXXXXXXXXXXXHQ, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, XXDXXXXXXXXXXXXXXXHV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXL, XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXQ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXH, XXDXXXXXXXXXXXXXXXXXXXXLXXQ, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXLQ, XXDXXXXXXXXXXYXXW, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHQ, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJL, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXLV, XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX, 
   XXDXXXXXXXXXXXXXXXXXL, XXDXXXXXXXXXXXXXXXXXXXXLXXV, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXP, XXDXXXXXXXXXXXXXXDDXXX, 
   XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXF, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXXLW, XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, 
   XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHL, XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
   XXDXXXXXXXXXXXXXWDXXXXXXXXXXXXXXXXXXX, XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXW, 
   XXDXXXXXXXXXXXXXXXXXXXXXXXFK, XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, 
   XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXV, XXDXXXXXXXXXXXXXXXXXXXXLXXW, 
   XXDXXXXXXXXXXYXXXK : std_logic;

begin
   caddr <= ( XXDDXXXXXX, XXDDXXXXXXF, XXDDXXXXX, XXDDXXXXXF, XXDDXXXXXH, 
      XXDDXXXXXJ, XXDDXXXXXK, XXDDXXXXXL, XXDDXXXXXP, XXDDXXXXXQ, XXDDXXXXXV, 
      XXDDXXXXXW );
   scrub_corrected <= XXXXXXXXXXXXXXDX;
   scrub_done <= XXXXXXDXXXX;
   
   XVXXX : VCC port map( Y => VXXXXXXXX);
   XYPXXXXX : BUFF port map( A => bypass, Y => XXYPXXXXXX);
   XXXXXXXXXX : AND2 port map( A => XXXXXXXXXLXXF, B => XXXDXXXXXXXXXXXXXXXXXX,
                           Y => correctable);
   XXXDX : GND port map( Y => XXDXXXXXX);
   XYPXXXXXF : BUFF port map( A => bypass, Y => XXYPXXXXXXF);
   XXXXXXXXXXF : AND2A port map( A => XXXXXXXXXLXXF, B => 
                           XXXDXXXXXXXXXXXXXXXXXX, Y => error);
   XYPXXXXXH : BUFF port map( A => bypass, Y => XXYPXXXXXXH);
   XXDXXXXXXXXXXXDXDXXXXXXXXXX : XOR2 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXFV, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXH, Y => XXDXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXDXDXXXXXXXX : XOR2 port map( A => wdata(17), B => wdata(8), Y 
                           => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXDXDXXXXXXXXF : XOR2 port map( A => wdata(6), B => wdata(4), Y 
                           => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXF : XOR4 port map( A => wdata(8), B => 
                           XXDXXXXXXXXXXXXXXXXXDXDX, C => wdata(19), D => 
                           wdata(13), Y => XXDXXXXXXXXXXXDXDXXXXXXXXFW);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXH : XOR2 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXHK, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXL, Y => XXDXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXDXDXXXXXXXXH : XOR2 port map( A => wdata(26), B => wdata(18), 
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXX : XOR4 port map( A => wdata(4), B => wdata(9),
                           C => XXDXXXXXXXXXXXDXDXXXXXXP, D => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXHF, Y => XXDXXXXXXXXXXXXXXL
                           );
   XXDXXXXXXXXXXXDXDXXXXXXXXXXJ : XOR4 port map( A => wdata(27), B => 
                           XXDXXXXXXXXXXXXXXXXXDXDX, C => wdata(12), D => 
                           wdata(17), Y => XXDXXXXXXXXXXXDXDXXXXXXXXHD);
   XXDXXXXXXXXXXXDXDXXXXXXXXJ : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXP, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX, C => wdata(15), D 
                           => wdata(18), Y => XXDXXXXXXXXXXXDXDXXXXXXJ);
   XXDXXXXXXXXXXXDXDXXXXXXXXK : XOR2 port map( A => wdata(25), B => wdata(21), 
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXK : CM8 port map( D0 => wdata(28), D1 => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXXXX, D3 => 
                           wdata(28), S00 => XXDXXXXXXXXXXXDXDXXXXXXJ, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXDXDXXXXXXXXHJ, S11 
                           => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXL : XOR4 port map( A => wdata(19), B => wdata(26)
                           , C => wdata(22), D => wdata(23), Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXHH);
   XXDXXXXXXXXXXXDXDXXXXXXXXL : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXW, B => wdata(12), C 
                           => wdata(7), D => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF, 
                           Y => XXDXXXXXXXXXXXDXDXXXXXXP);
   XXDXXXXXXXXXXXXXXDXD : XOR2 port map( A => wdata(2), B => wdata(0), Y => 
                           XXDXXXXXXXXXXXXXXXDXDX);
   XXDXXXXXXXXXXXDXDXXXXXXXXP : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXJ, B => wdata(12), C 
                           => wdata(5), D => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXP, 
                           Y => XXDXXXXXXXXXXXDXDXXXXXXF);
   XXDXXXXXXXXXXXDXDXXXXXXXXQ : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXK, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXH, C => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXFD, D => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXDXDXXXXXX);
   XXDXXXXXXXXXXXDXDXXXXXXXXV : XOR2 port map( A => wdata(23), B => wdata(13), 
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXDXDXXXXXXXXW : XOR2 port map( A => wdata(7), B => wdata(5), Y 
                           => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXDXDXXXXXXXXFD : XOR2 port map( A => wdata(16), B => wdata(11),
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXP : XOR4 port map( A => wdata(16), B => wdata(21)
                           , C => wdata(27), D => XXDXXXXXXXXXXXXXXXDXDX, Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXHF);
   XXDXXXXXXXXXXXDXDXXXXXXXXFF : XOR2 port map( A => wdata(22), B => wdata(20),
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXDXDXXXXXXXXFH : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXV, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXH, C => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXQ, D => wdata(19), Y 
                           => XXDXXXXXXXXXXXDXDXXXXXXL);
   XXDXXXXXXXXXXXDXDXXXXXXXXFJ : XOR2 port map( A => wdata(28), B => wdata(24),
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXDXDXXXXXXXXFK : XOR2 port map( A => wdata(15), B => wdata(10),
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXDXD : XOR2 port map( A => wdata(3), B => wdata(1), Y => 
                           XXDXXXXXXXXXXXXXXXXXDXDX);
   XXDXXXXXXXXXXXDXDXXXXXXXXFL : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXF, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXL, C => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXQ, D => wdata(6), Y 
                           => XXDXXXXXXXXXXXDXDXXXXXXK);
   XXDXXXXXXXXXXXDXDXXXXXXXXFP : XOR4 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXJ, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXX, C => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXW, D => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXV, Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXH);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXF : XOR4 port map( A => wdata(0), B => wdata(3)
                           , C => XXDXXXXXXXXXXXDXDXXXXXXF, D => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXHH, Y => XXDXXXXXXXXXXXXXX)
                           ;
   XXDXXXXXXXXXXXDXDXXXXXXXXFQ : XOR2 port map( A => wdata(14), B => wdata(9), 
                           Y => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXX : CM8INV port map( A => wdata(28), Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXQ : XOR2 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXHD, B => 
                           XXDXXXXXXXXXXXDXDXXXXXX, Y => XXDXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXV : XOR4 port map( A => wdata(10), B => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXFD, C => wdata(14), D
                           => XXDXXXXXXXXXXXXXXXDXDX, Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXHK);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXW : XOR2 port map( A => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXFW, B => 
                           XXDXXXXXXXXXXXDXDXXXXXXK, Y => XXDXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXFD : XOR4 port map( A => wdata(27), B => wdata(1)
                           , C => wdata(20), D => wdata(24), Y => 
                           XXDXXXXXXXXXXXDXDXXXXXXXXFV);
   XXDXXXXXXXXXXXDXDXXXXXXXXXXFF : XOR4 port map( A => wdata(11), B => 
                           wdata(25), C => XXDXXXXXXXXXXXDXDXXXXXXXXXXXXXXK, D 
                           => wdata(2), Y => XXDXXXXXXXXXXXDXDXXXXXXXXHJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => axrdata(12), Y =>
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXJF, D1 => 
                           XXDXXXXDXXXXXXXXH, D2 => XXDXXXXXX, D3 => VXXXXXXXX,
                           S00 => axrdata(29), S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S11 => 
                           XXDXXXXXXXX, Y => XXDXXXXXXXXXXKD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXHW, D1 
                           => XXDXXXXDXXXXXXXXK, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(3), S01 => VXXXXXXXX, S10 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S11
                           => XXDXXXXXXXXJ, Y => XXDXXXXXXXXXXJJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXHW, D1
                           => XXDXXXXDXXXXXXXXK, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(2), S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXH, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXJW);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => axrdata(23), Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D1 
                           => VXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S00
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX, S01 => VXXXXXXXX
                           , S10 => XXDXXXXDXXXXXYXXXXXXXXXXXXXH, S11 => 
                           XXDXXXXXX, Y => XXDXXXXDXXXXXXXXJ);
   XXDXXXXDXXXXXYXXXXXXX : XOR4 port map( A => axrdata(34), B => axrdata(27), C
                           => axrdata(30), D => axrdata(8), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => XXDXXXXXXXXXXV, 
                           Y => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXDXXXXXYXXXXXXXF : XOR2 port map( A => axrdata(16), B => axrdata(11), 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXFW);
   XXDXXXXDXXXXXYXXXXXXXH : XOR4 port map( A => axrdata(33), B => axrdata(26), 
                           C => axrdata(20), D => axrdata(10), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXV);
   XXDXXXXDXXXXXYXXXXXXXXX : XOR4 port map( A => axrdata(6), B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXL, C => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXP, D => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXQ, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : OR3A port map( A => 
                           XXDXXXXDXXXXXYXXXXXF, B => XXDXXXXDXXXXXYXXXXX, C =>
                           XXDXXXXDXXXXXYXXXXXJ, Y => XXDXXXXDXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXDXXXXXYXXXXXK, D1 => XXDXXXXXX, D2 => 
                           XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXDXXXXXYXXXXXK, S01 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXH, S11 => XXDXXXXXX, Y =>
                           XXDXXXXXXXXXXH);
   XXDXXXXDXXXXXYXXXXXXXXXF : XOR2 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXDXXXXXYXXXXXF);
   XXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXJ, Y => 
                           XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXH : AND3B port map( A => 
                           XXDXXXXDXXXXXYXXXXXF, B => XXDXXXXDXXXXXYXXXXXJ, C 
                           => XXDXXXXDXXXXXYXXXXX, Y => XXDXXXXXXXXXXV);
   XXDXXXXDXXXXXYXXXXXXXJ : XOR2 port map( A => axrdata(31), B => axrdata(24), 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => axrdata(27),
                           Y => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ)
                           ;
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXX : OR3B port map( A => XXDXXXXDXXXXXYXXXXXF, 
                           B => XXDXXXXDXXXXXYXXXXX, C => XXDXXXXDXXXXXXXXK, Y 
                           => XXDXXXXDXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXDXXXXXYXXXXXJ, 
                           D1 => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, D2 
                           => XXDXXXXXX, D3 => VXXXXXXXX, S00 => axrdata(34), 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXXXXJ, S11 => 
                           XXDXXXXDXXXXXXXXF, Y => XXDXXXXXXXXXXJH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => XXDXXXXXXXXXXFD, 
                           D1 => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW
                           , D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           axrdata(25), S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXXXXL, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXJD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXJF, 
                           D1 => XXDXXXXDXXXXXXXXH, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(16), S01 => VXXXXXXXX, S10
                           => XXDXXXXDXXXXXXXXL, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXFL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => axrdata(26)
                           , Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXXFLXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXDXXXXXXXFLXXXXXXXXXXXXXXXX, D1 => XXDXXXXXX, 
                           D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXDXXXXXXXFLXXXXXXXXXXXXXXXX, S01 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXH, S11 => XXDXXXXXX, Y =>
                           XXDXXXXXXXXXXHW);
   XXDXXXXDXXXXXYXXXXXXXXXXX : XOR4 port map( A => axrdata(17), B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXW, C => axrdata(12), D =>
                           axrdata(14), Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXFD, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8INV port map( A => axrdata(18)
                           , Y => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX
                           );
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => axrdata(12), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D2 => 
                           axrdata(12), D3 => axrdata(12), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXXXXXXXV, S10 => 
                           XXDXXXXDXXXXXYXXXXXXXHD, S11 => XXDXXXXDXXXXXXXXK, Y
                           => XXDXXXXXXXXXXK);
   XXDXXXXDXXXXXYXXXXXXXXXXXF : XOR4 port map( A => axrdata(24), B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFF, C => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXJ, D => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXK, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : OR2A port map( A => 
                           XXDXXXXDXXXXXYXXXXXF, B => XXDXXXXDXXXXXYXXXXX, Y =>
                           XXDXXXXDXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => axrdata(13), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D2 => 
                           axrdata(13), D3 => axrdata(13), S00 => 
                           XXDXXXXDXXXXXXXXXX, S01 => XXDXXXXXXXXXXFD, S10 => 
                           XXDXXXXDXXXXXYXXXXX, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXJK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => axrdata(20), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D2 => 
                           axrdata(20), D3 => axrdata(20), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXXXXXXXH, S10 => 
                           XXDXXXXDXXXXXXXX, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXW);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => axrdata(8), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, D2 => 
                           axrdata(8), D3 => axrdata(8), S00 => 
                           XXDXXXXDXXXXXYXXXXX, S01 => XXDXXXXDXXXXXXXXXX, S10 
                           => XXDXXXXDXXXXXXXXJ, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXHV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXL : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D2 
                           => VXXXXXXXX, D3 => XXDXXXXXXXXJ, S00 => 
                           XXDXXXXXXXXXXV, S01 => XXDXXXXXXXXXXFD, S10 => 
                           axrdata(22), S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXHQ)
                           ;
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXP : CM8 port map( D0 => XXDXXXXXXXXXXFD, 
                           D1 => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV
                           , D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           axrdata(32), S01 => VXXXXXXXX, S10 => XXDXXXXXXXXH, 
                           S11 => XXDXXXXXXXXF, Y => XXDXXXXXXXXXXHP);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXJ : XA1 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXH, C => 
                           XXDXXXXDXXXXXYXXXXXK, Y => XXDXXXXXXXXXXFD);
   XXDXXXXDXXXXXYXXXXXXXK : XOR2 port map( A => axrdata(33), B => axrdata(30), 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXFF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXF : OR2B port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXHD, B => XXDXXXXDXXXXXYXXXXXH, 
                           Y => XXDXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK : CM8INV port map( A => 
                           XXDXXXXXXXXJ, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXDXXXXXYXXXXXXXXXXXH : XOR4 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFV, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFH, C => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFL, D => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXDXXXXXYXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXL : CM8 port map( D0 => XXDXXXXXXXXXXH, D1 => 
                           XXDXXXXDXXXXXXXXJ, D2 => XXDXXXXXX, D3 => VXXXXXXXX,
                           S00 => axrdata(28), S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXXXXL, S11 => XXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXHK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXP : CM8 port map( D0 => axrdata(31), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D2 => 
                           axrdata(31), D3 => axrdata(31), S00 => 
                           XXDXXXXDXXXXXYXXXXX, S01 => XXDXXXXDXXXXXXXXXX, S10 
                           => XXDXXXXDXXXXXXXXK, S11 => XXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXFF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXQ : CM8 port map( D0 => axrdata(18), D1 =>
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D2 =>
                           axrdata(18), D3 => axrdata(18), S00 => 
                           XXDXXXXDXXXXXXXXXX, S01 => XXDXXXXXXXXXXJF, S10 => 
                           XXDXXXXDXXXXXYXXXXX, S11 => XXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXJQ);
   XXDXXXXDXXXXXYXXXXXXXXXH : XOR2 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXK, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFJ, Y => 
                           XXDXXXXDXXXXXYXXXXX);
   XXDXXXXDXXXXXYXXXXXXXL : XOR4 port map( A => XXDXXXXDXXXXXYXXXXXXXXXXXXXFF, 
                           B => XXDXXXXDXXXXXYXXXXXXXXXXXXXFQ, C => axrdata(34)
                           , D => axrdata(0), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXV : CM8INV port map( A => axrdata(15), Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXDXXXXXYXXXXXXXP : XOR2 port map( A => axrdata(12), B => axrdata(10), 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXW : CM8INV port map( A => XXDXXXXXXXXXXV, 
                           Y => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXYXXXXXXXQ : XOR2 port map( A => axrdata(35), B => axrdata(29), 
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXLXXXXXXXXXX : XOR2 port map( A => XXDXXXXDXXXXXYXXXXXH, 
                           B => XXDXXXXDXXXXXYXXXXXXXHD, Y => 
                           XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXX);
   XXDXXXXDXXXXXYXXXXXXXV : XOR2 port map( A => axrdata(17), B => axrdata(8), Y
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXFK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFD : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXJ, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXDXXXXXXFLXXXXXXXX : CM8 port map( D0 => XXDXXXXDXXXXXYXXXXXK, D1 => 
                           VXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXYXXXXXK, S00 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXDXXXXXYXXXXXXXXXXXXXH, S11 => 
                           XXDXXXXXX, Y => XXDXXXXDXXXXXXXXK);
   XXDXXXXDXXXXXYXXXXXXXW : XOR2 port map( A => axrdata(9), B => axrdata(7), Y 
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXW);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFF : CM8 port map( D0 => axrdata(30), D1 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, 
                           D2 => axrdata(30), D3 => axrdata(30), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXXXXXXXHW, S10 =>
                           XXDXXXXDXXXXXXXX, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXJF, D1
                           => XXDXXXXDXXXXXXXXH, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(6), S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXH, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXHL);
   XXDXXXXDXXXXXYXXXXXXXFD : XOR4 port map( A => axrdata(32), B => axrdata(28),
                           C => axrdata(23), D => axrdata(31), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFP);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => axrdata(5), 
                           Y => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXYXXXXXXXXXJ : XOR4 port map( A => axrdata(4), B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFH, C => axrdata(32), D 
                           => axrdata(22), Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXF)
                           ;
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFH : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXJ, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXK, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXLXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXF, Y => 
                           XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL : CM8INV port map( A => axrdata(11)
                           , Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFJ : CM8 port map( D0 => axrdata(26), D1 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, 
                           D2 => axrdata(26), D3 => axrdata(26), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXXXXXXXH, S10 => 
                           XXDXXXXDXXXXXYXXXXXXXHD, S11 => XXDXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXFJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXL : CM8INV port map( A => axrdata(8), Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH);
   XXDXXXXDXXXXXYXXXXXXXFF : XOR2 port map( A => axrdata(23), B => axrdata(20),
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXFV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXQ : CM8 port map( D0 => XXDXXXXXXXXXXH, D1 => 
                           XXDXXXXDXXXXXXXXJ, D2 => XXDXXXXXX, D3 => VXXXXXXXX,
                           S00 => axrdata(33), S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXXXXL, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXFH);
   XXDXXXXDXXXXXYXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFK : CM8 port map( D0 => XXDXXXXXXXXXXJF, 
                           D1 => XXDXXXXDXXXXXXXXH, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(35), S01 => VXXXXXXXX, S10
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, 
                           S11 => XXDXXXXXXXXF, Y => XXDXXXXXXXXXXHH);
   XXDXXXXDXXXXXYXXXXXXXXXK : XOR4 port map( A => XXDXXXXDXXXXXYXXXXXXXXXXXXXFK
                           , B => XXDXXXXDXXXXXYXXXXXXXXXXXXXP, C => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXHD, D => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXJ, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFL : CM8 port map( D0 => axrdata(27), D1 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, 
                           D2 => axrdata(27), D3 => axrdata(27), S00 => 
                           XXDXXXXDXXXXXYXXXXX, S01 => XXDXXXXDXXXXXXXXXX, S10 
                           => XXDXXXXDXXXXXXXXH, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXHD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFP : CM8 port map( D0 => axrdata(11), D1 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, 
                           D2 => axrdata(11), D3 => axrdata(11), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXXXXXXXJF, S10 =>
                           XXDXXXXDXXXXXXXX, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXP);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXV : CM8 port map( D0 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D1 => 
                           XXDXXXXDXXXXXYXXXXXJ, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(19), S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXX, S11 => XXDXXXXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXX);
   XXDXXXXDXXXXXYXXXXXXXXXXXJ : XOR2 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXJ, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFW, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP : CM8INV port map( A => axrdata(21)
                           , Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXP : CM8 port map( D0 => axrdata(5), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D2 =>
                           axrdata(5), D3 => axrdata(5), S00 => 
                           XXDXXXXDXXXXXXXXXX, S01 => XXDXXXXXXXXXXHW, S10 => 
                           XXDXXXXDXXXXXYXXXXX, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXHF);
   XXDXXXXDXXXXXYXXXXXXXFH : XOR4 port map( A => axrdata(26), B => axrdata(7), 
                           C => axrdata(2), D => axrdata(19), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => VXXXXXXXX, D1 =>
                           XXDXXXXDXXXXXYXXXXXK, D2 => XXDXXXXDXXXXXYXXXXXK, D3
                           => VXXXXXXXX, S00 => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX
                           , S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXH, S11 => XXDXXXXXX, Y =>
                           XXDXXXXDXXXXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXV, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXQ : CM8INV port map( A => axrdata(7), Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ);
   XXDXXXXDXXXXXYXXXXXXXXXL : XOR4 port map( A => axrdata(35), B => axrdata(1),
                           C => XXDXXXXDXXXXXYXXXXXXXXXXXXXQ, D => axrdata(26),
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => XXDXXXXXX, D1 
                           => VXXXXXXXX, D2 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
                           D3 => XXDXXXXXX, S00 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, 
                           S01 => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXH, S11 => XXDXXXXXX, Y =>
                           XXDXXXXXXXXXXJF);
   XXDXXXXDXXXXXYXXXXXXXFJ : XOR4 port map( A => XXDXXXXDXXXXXYXXXXXXXXXXXXXF, 
                           B => XXDXXXXDXXXXXYXXXXXXXXXXXXXL, C => axrdata(34),
                           D => axrdata(3), Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXFJ)
                           ;
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXV : CM8 port map( D0 => XXDXXXXXXXXXXH, D1 
                           => XXDXXXXDXXXXXXXXJ, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(4), S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXH, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXJV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFQ : CM8INV port map( A => axrdata(31), Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXDXXXXXYXXXXXXXFK : XOR2 port map( A => axrdata(28), B => axrdata(25),
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXFQ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXW : CM8 port map( D0 => XXDXXXXXXXXXXJF, D1
                           => XXDXXXXDXXXXXXXXH, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(9), S01 => VXXXXXXXX, S10 
                           => XXDXXXXDXXXXXXXXL, S11 => XXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXFV);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXFD : CM8 port map( D0 => XXDXXXXXXXXXXHW, 
                           D1 => XXDXXXXDXXXXXXXXK, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(0), S01 => VXXXXXXXX, S10 
                           => XXDXXXXDXXXXXXXXL, S11 => XXDXXXXXXXXJ, Y => 
                           XXDXXXXXXXXXXJP);
   XXDXXXXDXXXXXYXXXXXXXXXXXK : XOR4 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFQ, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFK, C => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXV, D => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXDXXXXXYXXXXXK);
   XXDXXXXDXXXXXXXXXXXXLXXXXXX : CM8 port map( D0 => 
                           XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXX, D1 => 
                           XXDXXXXDXXXXXYXXXXXF, D2 => XXDXXXXDXXXXXYXXXXXF, D3
                           => XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXX, S00 => 
                           XXDXXXXDXXXXXXXXXXF, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXYXXXXX, S11 => XXDXXXXXX, Y => 
                           XXXXXXXXXLXXF);
   XXDXXXXDXXXXXXFLXXXXXXXXXXXXXXX : CM8INV port map( A => XXDXXXXDXXXXXYXXXXXK
                           , Y => XXDXXXXDXXXXXXXFLXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXW : CM8 port map( D0 => axrdata(15), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, D2 => 
                           axrdata(15), D3 => axrdata(15), S00 => 
                           XXDXXXXDXXXXXXXXXX, S01 => XXDXXXXXXXXXXH, S10 => 
                           XXDXXXXDXXXXXYXXXXX, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXFK);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFV : CM8 port map( D0 => axrdata(24), D1 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, 
                           D2 => axrdata(24), D3 => axrdata(24), S00 => 
                           XXDXXXXDXXXXXYXXXXX, S01 => XXDXXXXDXXXXXXXXXX, S10 
                           => XXDXXXXDXXXXXXXXK, S11 => XXDXXXXXXXX, Y => 
                           XXDXXXXXXXXXXJL);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXFW : CM8 port map( D0 => XXDXXXXXXXXXXH, 
                           D1 => XXDXXXXDXXXXXXXXJ, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(17), S01 => VXXXXXXXX, S10
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, 
                           S11 => XXDXXXXXXXXF, Y => XXDXXXXXXXXXXFQ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXFF : AND2A port map( A => 
                           XXDXXXXDXXXXXYXXXXXF, B => XXDXXXXDXXXXXYXXXXXJ, Y 
                           => XXDXXXXDXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXFD : CM8 port map( D0 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, D1 => 
                           XXDXXXXDXXXXXYXXXXXJ, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(14), S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXXF, S11 => XXDXXXXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXF);
   XXDXXXXDXXXXXYXXXXXXXXXXXXX : XNOR2 port map( A => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXX, Y => 
                           XXDXXXXDXXXXXYXXXXXXXHD);
   XXDXXXXDXXXXXYXXXXXXXFL : XOR2 port map( A => axrdata(19), B => axrdata(14),
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXHD);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXK : OR2 port map( A => 
                           XXDXXXXDXXXXXYXXXXXH, B => XXDXXXXDXXXXXYXXXXXXXHD, 
                           Y => XXDXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXHD : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXJ, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXDXXXXXYXXXXXXXFP : XOR2 port map( A => axrdata(21), B => axrdata(18),
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXQ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXHF : CM8INV port map( A => axrdata(20), Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXDXXXXXYXXXXXXXFQ : XOR4 port map( A => axrdata(32), B => axrdata(13),
                           C => axrdata(25), D => axrdata(9), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXHH : CM8INV port map( A => axrdata(13), Y 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXYXXXXXXXFV : XOR2 port map( A => axrdata(15), B => axrdata(13),
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXFH);
   XXDXXXXDXXXXXYXXXXXXXFW : XOR2 port map( A => axrdata(27), B => axrdata(22),
                           Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXP);
   XXDXXXXDXXXXXYXXXXXXXXXP : XOR4 port map( A => axrdata(5), B => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXF, C => axrdata(11), D =>
                           axrdata(18), Y => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXP);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXFH : CM8 port map( D0 => XXDXXXXXXXXXXHW, 
                           D1 => XXDXXXXDXXXXXXXXK, D2 => XXDXXXXXX, D3 => 
                           VXXXXXXXX, S00 => axrdata(1), S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXH, S11 => XXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXQ);
   XXDXXXXDXXXXXXFLXXXXXX : OR2A port map( A => XXDXXXXDXXXXXYXXXXXXXHD, B => 
                           XXDXXXXDXXXXXYXXXXXH, Y => XXDXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => axrdata(7), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, D2 => 
                           axrdata(7), D3 => axrdata(7), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXXXXXXXHW, S10 =>
                           XXDXXXXDXXXXXYXXXXXXXHD, S11 => XXDXXXXDXXXXXXXXL, Y
                           => XXDXXXXXXXXXXJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV : CM8INV port map( A => axrdata(30)
                           , Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXHJ : CM8 port map( D0 => axrdata(21), D1 
                           => XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, 
                           D2 => axrdata(21), D3 => axrdata(21), S00 => 
                           XXDXXXXDXXXXXYXXXXXH, S01 => XXDXXXXXXXXXXJF, S10 =>
                           XXDXXXXDXXXXXYXXXXXXXHD, S11 => XXDXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXFW);
   XXDXXXXDXXXXXYXXXXXXXXXXXL : CM8 port map( D0 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXF, D1 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXXXXXX, D3 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXXXF, S00 => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFP, S01 => VXXXXXXXX, S10
                           => XXDXXXXDXXXXXYXXXXXXXXXXXXXXXL, S11 => XXDXXXXXX,
                           Y => XXDXXXXDXXXXXYXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXDXXXXXYXXXXXK, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW : CM8INV port map( A => 
                           XXDXXXXXXXXXXV, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXDXXXXXXFLXXXXXXXXF : OR3 port map( A => XXDXXXXDXXXXXYXXXXX, B => 
                           XXDXXXXDXXXXXYXXXXXF, C => XXDXXXXDXXXXXYXXXXXJ, Y 
                           => XXDXXXXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD : CM8INV port map( A => 
                           axrdata(24), Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXDXXXXXXXXXXXXLXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXXXX, D1 => 
                           XXDXXXXDXXXXXYXXXXXJ, D2 => XXDXXXXDXXXXXYXXXXXJ, D3
                           => XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXXXXX, S00 => 
                           XXDXXXXDXXXXXXXXXXXXXLXXXXXXXXXXX, S01 => VXXXXXXXX,
                           S10 => XXDXXXXXXXXXXFD, S11 => XXDXXXXXXXXXXHW, Y =>
                           XXDXXXXDXXXXXXXXXXF);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXFF : CM8 port map( D0 => axrdata(23), D1 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, D2 => 
                           axrdata(23), D3 => axrdata(23), S00 => 
                           XXDXXXXDXXXXXYXXXXXJ, S01 => XXDXXXXXXXXXXHW, S10 =>
                           XXDXXXXDXXXXXXXX, S11 => XXDXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXFP);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXFH : CM8 port map( D0 => XXDXXXXXXXXXXH, D1 => 
                           XXDXXXXDXXXXXXXXJ, D2 => XXDXXXXXX, D3 => VXXXXXXXX,
                           S00 => axrdata(10), S01 => VXXXXXXXX, S10 => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, S11 => 
                           XXDXXXXXXXX, Y => XXDXXXXXXXXXXHJ);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXV, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXDXXXXXYXXXXXXXXXQ : XOR4 port map( A => XXDXXXXDXXXXXYXXXXXXXXXXXXXHD
                           , B => XXDXXXXDXXXXXYXXXXXXXXXXXXXFV, C => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXW, D => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXFW, Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXXH);
   XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF : CM8INV port map( A => 
                           XXDXXXXXXXXXXFD, Y => 
                           XXDXXXXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXDXXXXXYXXXXXXXXXV : XOR4 port map( A => axrdata(29), B => axrdata(16)
                           , C => axrdata(21), D => axrdata(15), Y => 
                           XXDXXXXDXXXXXYXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXXXXXXXX : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHD, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF);
   XXDXXXXXXXXXXXXXXXXXXXXX : OR2 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => rds(2), Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXWDXXXXXXXX : DFE3C port map( D => XXDXXXXXXXXXXFL, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXWDXXXXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXJD, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => XXXXXXXXXLXXF, D1 => 
                           VXXXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S11 
                           => XXDXXXXXXXXXXXXXXXW, Y => XXDXXXXXXXXXXYXXXF);
   XXDXXXXXXXXXXXXXXXXXXXLXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKL, D1 => tmout(19), D2 
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S01 => VXXXXXXXX,
                           S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFK);
   XXDXXXXXXXXXXXXXDDXXLX : XA1 port map( A => XXDDXXXXXW, B => XXDDXXXXXV, C 
                           => XXDXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXP);
   XXDXXXXXXXXXXXXXXXXXXXLXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFK, D1 => tmout(30),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, D3 => 
                           tmout(30), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXK);
   XXDXXXXXXXXXXXXXWDXXXXXXXX : CM8 port map( D0 => wdata(20), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXW, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(27));
   XXDXXXXXXXXXXXXWDXXXXXXXXH : DFE3C port map( D => XXDXXXXXXXXXXFQ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFH);
   XXDXXXXXXXXXXXXDXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXHV, D1 => 
                           axrdata(8), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rdata(1));
   XXDXXXXXXXXXXXXXXXXXXXLXXH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH, D2 => tmout(17), D3 
                           => tmout(17), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => XXDXXXXXX,
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXP);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFD, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXWDXXXXXXXXJ : DFE3C port map( D => XXDXXXXXXXXXXJL, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFV);
   XXDXXXXXXXXXXXXDXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXJ, D1 => 
                           axrdata(7), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rdata(0));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXP);
   XXDXXXXXXXXXXXXXWDXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXXXXXH, D1 => 
                           wp(6), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXK, D3 => 
                           XXDXXXXXX, S00 => XXYPXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S11 => XXDXXXXXX, Y 
                           => axwdata(6));
   XXDXXXXXXXXXXXXXWXDDXXXXX : CM8 port map( D0 => waddr(4), D1 => XXDDXXXXXL, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(4));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXH : AND4B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXL, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXXXXX : OR4A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKF);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXF, D1 
                           => XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXF, S00 
                           => XXDDXXXXXJ, S01 => VXXXXXXXX, S10 => waddr(6), 
                           S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXL);
   XXDXXXXXXXXXXXXXXDDXXXXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXV, E
                           => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn, Q
                           => XXDDXXXXXH);
   XXDXXXXXXXXXXXXXXXDDXXXXXX : CM8 port map( D0 => raddr(11), D1 => XXDDXXXXXX
                           , D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(11));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXX : CM8 port map( D0 => axrdata(35), D1 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXH, D2 => 
                           axrdata(35), D3 => axrdata(35), S00 => 
                           XXDXXXXXXXXXXV, S01 => XXDXXXXXXXXXXJF, S10 => 
                           XXYPXXXXXXF, S11 => XXDXXXXXXXXF, Y => rdata(28));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8INV port map( A => XXDXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXDDXX : AND2A port map( A => bypass, B => 
                           XXDXXXXXXXXXXXXXXXHK, Y => XXDXXXXXXXXXXXXXXDDXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, D2 => XXDXXXXXX
                           , D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJL, S01 => 
                           VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLD);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXX : CM8INV port map( A => axrdata(29), Y =>
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXXF : CM8 port map( D0 => wdata(7), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFH, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(14));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXX : OR2A port map( A => XXDXXXXXXXXXXYXXQ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXYXXXJ);
   XXDXXXXXXXXXXXXXDDXXLXF : AND2 port map( A => XXDXXXXXXXXXXXXXXXXXH, B => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXX : AND2A port map( A => 
                           XXDXXXXXXXXXXYXXV, B => XXXXXXDXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXP, D1 => tmout(39), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, D3 => 
                           tmout(39), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXH);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => axrdata(17), Y 
                           => XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXQ, D1 => tmout(22), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, D3 => 
                           tmout(22), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFP);
   XXDXXXXXXXXXXXXXWDXXXXXXXXH : CM8 port map( D0 => wdata(19), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHK, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(26));
   XXDXXXXXXXXXXXXXDDXXXXX : AND4 port map( A => XXDDXXXXXL, B => XXDDXXXXXK, C
                           => XXDDXXXXXJ, D => XXDDXXXXXH, Y => 
                           XXDXXXXXXXXXXYXXXH);
   XXDXXXXXXXXXXXXXWDXXXXXXXXJ : CM8 port map( D0 => wdata(8), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHD, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(15));
   XXDXXXXXXXXXXXXXXDDXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXF, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXJ);
   XXDXXXXXXXXXXXXXWXDDXXXXXF : CM8 port map( D0 => waddr(5), D1 => XXDDXXXXXK,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(5));
   XXDXXXXXXXXXXXXXXXDDXXXXXXF : CM8 port map( D0 => raddr(10), D1 => 
                           XXDDXXXXXXF, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10
                           => XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(10));
   XXDXXXXXXXXXXXXXXXXXXXXXXH : OR4 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKK, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJW);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXLX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXL, D1 => tmout(6), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, D3 => 
                           tmout(6), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 
                           => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXFF, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXJ);
   XXDXXXXXXXXXXXXXWDXXXXXXXF : CM8 port map( D0 => wdata(0), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXV, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(7));
   XXDXXXXXXXXXXXXXWDXXXXXXXXK : CM8 port map( D0 => wdata(25), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXV, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(32));
   XXDXXXXXXXXXXXXXXXXXXXX : AND2A port map( A => XXDXXXXXXXXXXYXXV, B => 
                           XXDXXXXXXXXXXYXX, Y => XXDXXXXXXXXXXXXXXXHQ);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXX : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXX, S01 => 
                           XXDXXXXXXXXXXYXXJ, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX, S11 => 
                           XXDXXXXXXXXXXXXXXXFJ, Y => XXDXXXXXXXXXXYXXH);
   XXDXXXXXXXXXXXXXWDXXXXXXXXL : CM8 port map( D0 => wdata(11), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHL, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(18));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXH : OR4A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXXXXXXXXJ : OR4 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLP, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJL, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, D1 => XXDXXXXXX
                           , D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, S01 => VXXXXXXXX
                           , S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, S11 =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXV, D1 => tmout(1), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D3 => tmout(1)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ
                           , S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXW
                           );
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXL : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHL);
   XXDXXXXXXXXXXXXXWXDDXXXXXH : CM8 port map( D0 => waddr(8), D1 => XXDDXXXXXF,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(8));
   XXDXXXXXXXXXXXXXXX : XOR2 port map( A => XXDDXXXXX, B => waddr(9), Y => 
                           XXDXXXXXXXXXXXXXXXHD);
   XXDXXXXXXXXXXXXXDDXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXXXXXX, D2 => VXXXXXXXX, D3 
                           => XXDXXXXXXXXXXYXXXK, S00 => XXDDXXXXXL, S01 => 
                           XXDDXXXXXK, S10 => XXDDXXXXXJ, S11 => XXDXXXXXX, Y 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXLXXL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFD, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, D2 => tmout(25)
                           , D3 => tmout(25), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKJ, S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHK);
   XXDXXXXXXXXXXXXXXWXXXXXXXX : AND2B port map( A => re, B => we, Y => 
                           XXDXXXXXXXXXXXXXXXHK);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXFF, D1 => 
                           axrdata(31), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXF, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(24));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXJL, D1 => 
                           axrdata(24), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(17));
   XXDXXXXXXXXXXXXXDDXLDXXXXXXXX : AND3B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLK, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLV, C => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXYXXW);
   XXDXXXXXXXXXXXXXXXDDXXXXX : CM8 port map( D0 => raddr(2), D1 => XXDDXXXXXQ, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(2));
   XXDXXXXXXXXXXXXWDXXXXXXX : DFE3C port map( D => XXDXXXXXXXXXXJW, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXWDXXXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXJJ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXX, D1 => VXXXXXXXX, D2
                           => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXHL, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLV, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJF, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJL);
   XXDXXXXXXXXXXXXPXXXXXXXXX : CM8INV port map( A => axrdata(3), Y => 
                           XXDXXXXXXXXXXXXPXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWXDDXXXXXJ : CM8 port map( D0 => waddr(9), D1 => XXDDXXXXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(9));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXYXX, 
                           D1 => VXXXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX,
                           S01 => XXDXXXXXXXXXXXXXXXFQ, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX : AND3 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXQXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXX, E => XXDXXXXXXXXXXYXXK,
                           CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXDDXXXXXF : CM8 port map( D0 => raddr(3), D1 => XXDDXXXXXP,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(3));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXJ : CM8 port map( D0 => XXDXXXXXXXXXXHP, D1 => 
                           axrdata(32), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXF, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(25));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXV : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXFP, D1 => 
                           axrdata(23), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(16));
   XXDXXXXXXXXXXXXXWDXXXXXXXXP : CM8 port map( D0 => wdata(12), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXQ, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(19));
   XXDXXXXXXXXXXXXXDDXXXXF : AND2A port map( A => XXYPXXXXXXF, B => 
                           XXDXXXXXXXXXXXXXXXHK, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFL);
   XXDXXXXXXXXXXXXXDDXXLXH : XA1 port map( A => XXDXXXXXXXXXXXXXXXFF, B => 
                           XXDDXXXXXF, C => XXDXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXL);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXW : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXX : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXK, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV);
   XXDXXXXXXXXXXXXXWDXXXXXXXXQ : CM8 port map( D0 => wdata(26), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHH, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(33));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFD : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFP, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFL, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH);
   XXDXXXXXXXXXXXXXXXXXXXLXH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, D1 => tmout(8), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, D3 => tmout(8)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF,
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXV);
   XXDXXXXXXXXXXXXXXXXXXXXF : AND2B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, B => 
                           XXDXXXXXXXXXXYXXV, Y => XXDXXXXXXXXXXXXXXXHF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXL, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXWDXXXXXXXXK : DFE3C port map( D => XXDXXXXXXXXXXHK, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXPXXXX : CM8 port map( D0 => XXDXXXXXXXXXXJW, D1 => axrdata(2)
                           , D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => bypass, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => rp(2));
   XXDXXXXXXXXXXXXXXXF : XOR2 port map( A => XXDDXXXXXW, B => waddr(0), Y => 
                           XXDXXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXK);
   XXDXXXXXXXXXXXXWDXXXXXXXXL : DFE3C port map( D => XXDXXXXXXXXXXKD, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFW);
   XXDXXXXXXXXXXXXWDXXXXXXXXP : DFE3C port map( D => XXDXXXXXXXXXXL, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, D2 => XXDXXXXXX,
                           D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, S01 => 
                           VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLQ);
   XXDXXXXXXXXXXXXWDXXXXXXXXQ : DFE3C port map( D => XXDXXXXXXXXXXFF, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXL, D1 => tmout(10), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, D3 => 
                           tmout(10), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01
                           => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXFK, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFV
                           );
   XXDXXXXXXXXXXXXPXXXXF : CM8 port map( D0 => axrdata(3), D1 => 
                           XXDXXXXXXXXXXXXPXXXXXXXXXXXXXXX, D2 => axrdata(3), 
                           D3 => axrdata(3), S00 => XXDXXXXXXXXXXV, S01 => 
                           XXDXXXXXXXXXXHW, S10 => bypass, S11 => XXDXXXXXXXXJ,
                           Y => rp(3));
   XXDXXXXXXXXXXXXXXXXXXXLXXQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXJ, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, D2 => tmout(37)
                           , D3 => tmout(37), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKQ, S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHD);
   XXDXXXXXXXXXXXXXXWXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXHD, D1 => 
                           VXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXHD, S00 => XXDDXXXXXX, S01 => 
                           VXXXXXXXX, S10 => waddr(11), S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFW, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFD : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFV, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXW);
   XXDXXXXXXXXXXXXXWXDDXXXXXK : CM8 port map( D0 => waddr(0), D1 => XXDDXXXXXW,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(0));
   XXDXXXXXXXXXXXXXWXDDXXXXXL : CM8 port map( D0 => waddr(1), D1 => XXDDXXXXXV,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(1));
   XXDXXXXXXXXXXXXXXXH : XOR2 port map( A => XXDDXXXXXF, B => waddr(8), Y => 
                           XXDXXXXXXXXXXXXXXXFV);
   XXDXXXXXXXXXXXXXXXXXXXLXXV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, D1 => tmout(18)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXW, D3 => 
                           tmout(18), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH, S11 => XXDXXXXXX, Y 
                           => XXDXXXXXXXXXXXXXXXXXXXXLXXXFH);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXDDXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXL : OR4A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKH);
   XXDXXXXXXXXXXXXXDDXXXXH : AND2A port map( A => XXYPXXXXXXF, B => 
                           XXDXXXXXXXXXXXXXXXHK, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFD);
   XXDXXXXXXXXXXXXXWDXXXXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXXXXXF, D1 => 
                           wp(3), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXW, D3 => 
                           XXDXXXXXX, S00 => XXYPXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S11 => XXDXXXXXX, Y 
                           => axwdata(3));
   XXDXXXXXXXXXXXXXXXXXXXXXXP : OR3 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKV, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKD);
   XXDXXXXXXXXXXXXXXDDXXXXXH : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXX, E
                           => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn, Q
                           => XXDDXXXXXQ);
   XXDXXXXXXXXXXXXXWDXXXXXXXXV : CM8 port map( D0 => wdata(15), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHF, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(22));
   XXDXXXXXXXXXXXXXWDXXXXXXXXW : CM8 port map( D0 => wdata(4), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHJ, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(11));
   XXDXXXXXXXXXXFXXXXLXXD : DFP1B port map( D => XXDXXXXXX, CLK => clk, PRE => 
                           rstn, Q => XXDXXXXXXXXXXXFXXXXLXXDX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXDDXLDXXXXXXXXXX : AND2 port map( A => XXDXXXXXXXXXXYXX, B =>
                           XXDXXXXXXXXXXXXXXXDDXX, Y => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXXLXXW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFH, D1 => tmout(24),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, D3 => 
                           tmout(24), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXQ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => axrdata(22), Y 
                           => XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => XXDXXXXXX, D2 
                           => VXXXXXXXX, D3 => XXDXXXXXXXXJ, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXF, S01 => 
                           XXDXXXXXXXXXXHW, S10 => stop_scrub, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXXDXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXXFD : CM8 port map( D0 => wdata(16), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFF, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(23));
   XXDXXXXXXXXXXXXXWDXXXXXXXXFF : CM8 port map( D0 => wdata(3), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFD, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(10));
   XXDXXXXXXXXXXXXXDDXXLXJ : AND2A port map( A => XXDDXXXXXW, B => 
                           XXDXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXDDXXXXJ : AND2A port map( A => XXDXXXXXXXXXXYXXXK, B => 
                           XXDXXXXXXXXXXYXXXH, Y => XXDXXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXXDDXXLXXXXXX : CM8INV port map( A => XXDDXXXXXJ, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXFD : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXV, D1 => tmout(31), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, D3 => 
                           tmout(31), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXJW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHW);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXK, D1 => 
                           axrdata(12), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(5));
   XXDXXXXXXXXXXXXXXXXXXXLXJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXQ, D1 => tmout(0), D2
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => VXXXXXXXX, S10
                           => XXDXXXXXX, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXF);
   XXDXXXXXXXXXXXXXDDXXLXK : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXH, D2 => XXDXXXXXXXXXXXXXXXXXH, 
                           D3 => XXDXXXXXX, S00 => XXDDXXXXXF, S01 => 
                           XXDXXXXXXXXXXXXXXXFF, S10 => XXDDXXXXX, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXDDXXLXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFF : AND3B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXWDXXXXXXXJ : CM8 port map( D0 => XXDXXXXXXXXXXXXXX, D1 => 
                           wp(2), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXJ, D3 => 
                           XXDXXXXXX, S00 => XXYPXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S11 => XXDXXXXXX, Y 
                           => axwdata(2));
   XXDXXXXXXXXXXXXXXDDXXXXXJ : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXW, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXP);
   XXDXXXXXXXXXXXXWDXXXXXXXXV : DFE3C port map( D => XXDXXXXXXXXXXJK, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFQ);
   XXDXXXXXXXXXXXXWDXXXXXXXXW : DFE3C port map( D => XXDXXXXXXXXXXW, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXLXXFF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXF, D1 => tmout(11), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, D3 => 
                           tmout(11), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01
                           => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFH, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXF : AND4C port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFD, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXQ : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXFL, D1 =>
                           VXXXXXXXX, D2 => VXXXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXFL, S00 => XXDDXXXXXX, S01 => 
                           VXXXXXXXX, S10 => rds(3), S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFJ, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXFH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXK, D1 => tmout(36), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, D3 => 
                           tmout(36), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFD);
   XXDXXXXXXXXXXXXDXXXXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXP, D1 => 
                           axrdata(11), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(4));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFQ, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX : AND2B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXYXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHF, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXP, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : OR2B port map( A => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFD, B => 
                           XXDXXXXXXXXXXXXXXXFH, Y => XXDXXXXXXXXXXXXXXXFQ);
   XXDXXXXXXXXXXXXWDXXXXXXXXFD : DFE3C port map( D => XXDXXXXXXXXXXK, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFK, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXXJ : XOR2 port map( A => XXDDXXXXXV, B => waddr(1), Y => 
                           XXDXXXXXXXXXXXXXXXHP);
   XXDXXXXXXXXXXXXLXWDXWXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXXFLXX, E => 
                           XXDXXXXXXXXXXYXXV, CLK => clk, CLR => rstn, Q => 
                           slowdown);
   XXDXXXXXXXXXXXXWDXXXXXXXXFF : DFE3C port map( D => XXDXXXXXXXXXXFW, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXWXXXXX : CM8 port map( D0 => waddr(10), D1 => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXXXXX, D2 => VXXXXXXXX, D3 
                           => VXXXXXXXX, S00 => XXDDXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXXFV, S11 => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXX, Y => XXDXXXXXXXXXXY);
   XXDXXXXXXXXXXXXXXXXXXXXXXV : OR3 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKJ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKK);
   XXDXXXXXXXXXXXXXXXXXXXLXK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXK, D1 => tmout(9), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, D3 => 
                           tmout(9), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 
                           => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXX);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXX, D1 =>
                           waddr(7), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDDXXXXXH, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXHP, S11 => XXDXXXXXXXXXXXXXXXHH, Y
                           => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, S01 => 
                           VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP);
   XXDXXXXXXXXXXXXXDDXXXXXXXXX : OR2B port map( A => XXDDXXXXXV, B => 
                           XXDDXXXXXW, Y => XXDXXXXXXXXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHH, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, S01 => 
                           VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXYXXQ, 
                           D1 => VXXXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, S11 => 
                           XXDXXXXXXXXXXXXXXXXXF, Y => XXDXXXXXXXXXXYXXP);
   XXDXXXXXXXXXXXXWDXXXXXXXXFH : DFE3C port map( D => XXDXXXXXXXXXXHH, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXH : AND3B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXWDXXXXXXXXFJ : DFE3C port map( D => XXDXXXXXXXXXXJH, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXXXXXXXXLK,
                           D1 => VXXXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXLV, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXYXXV, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXPXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXHL, D1 => 
                           axrdata(6), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rp(6));
   XXDXXXXXXXXXXXXXDDXXXXK : AND4A port map( A => XXDXXXXXXXXXXYXXXK, B => 
                           XXDDXXXXX, C => XXDXXXXXXXXXXYXXXH, D => XXDDXXXXXF,
                           Y => XXDXXXXXXXXXXXXXXDDXXXXXFJ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXL : CM8 port map( D0 => XXDXXXXXXXXXXW, D1 => 
                           axrdata(20), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(13));
   XXDXXXXXXXXXXXXXXXXXXXXXF : OR4A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFJ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXJ, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXXXLXXFJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, D1 => tmout(16)
                           , D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFJ, D3 => 
                           tmout(16), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, S11 => XXDXXXXXX, 
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFF, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK);
   XXDXXXXXXXXXXXXXDDXXLXL : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXH, S00 => XXDDXXXXXH, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXDDXXLXXXXXXX, S11
                           => XXDXXXXXXXXXXXXXXDDXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXV);
   XXDXXXXXXXXXXXXXXXXXXXLXL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXP, D1 => tmout(7), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D3 => 
                           tmout(7), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 
                           => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXP);
   XXDXXXXXXXXXXXXXXXXXXXXXH : DFC1B port map( D => XXDXXXXXXXXXXYXXXF, CLK => 
                           clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXFW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXW, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHD : AND3B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXW : OR3 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKK, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLW);
   XXDXXXXXXXXXXXXXXXDDXXXXXH : CM8 port map( D0 => raddr(7), D1 => XXDDXXXXXH,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(7));
   XXDXXXXXXXXXXXXXXXXDXXXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXXHF, E => 
                           XXDXXXXXXXXXXYXXP, CLK => clk, CLR => rstn, Q => 
                           XXXXXXDXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXFK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXH, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, D2 => tmout(23),
                           D3 => tmout(23), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKW, S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFW);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXP : CM8 port map( D0 => XXDXXXXXXXXXXHK, D1 => 
                           axrdata(28), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXF, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(21));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXF : CM8 port map( D0 => XXDXXXXXXXXXXFK, D1 => 
                           axrdata(15), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(8));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXQ : CM8 port map( D0 => XXDXXXXXXXXXX, D1 => 
                           axrdata(19), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(12));
   XXDXXXXXXXXXXXXWDXXXXXXXH : DFE3C port map( D => XXDXXXXXXXXXXHL, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXWX : DFC1B port map( D => XXDXXXXXXXXXXYXXF, CLK => clk, CLR 
                           => rstn, Q => XXDXXXXXXXXXXXXWXX);
   XXDXXXXXXXXXXXXWDXXXXXXXJ : DFE3C port map( D => XXDXXXXXXXXXXJ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXXXDDXXXXXJ : CM8 port map( D0 => raddr(6), D1 => XXDDXXXXXJ,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(6));
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXX : OR3A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, B => 
                           XXDXXXXXXXXXXYXXV, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXV : CM8 port map( D0 => XXDXXXXXXXXXXHD, D1 => 
                           axrdata(27), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXF, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(20));
   XXDXXXXXXXXXXXXXXXXXXXLXXFL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXX, D1 => tmout(38), 
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, D3 => 
                           tmout(38), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHP);
   XXDXXXXXXXXXXXXXXXXXXXXXJ : DFC1B port map( D => XXDXXXXXXXXXXYXXX, CLK => 
                           clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXH : CM8 port map( D0 => XXDXXXXXXXXXXFL, D1 => 
                           axrdata(16), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(9));
   XXDXXXXXXXXXXXXXXXXXXXXXXFD : OR3A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLH);
   XXDXXXXXXXXXXXXXWDXXXXXXXXXXXXX : CM8INV port map( A => XXDXXXXXXXXXXXXXXXHK
                           , Y => XXDXXXXXXXXXXXXXWDXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHH);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX, D2 => 
                           XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXH, S10 => 
                           XXDXXXXXXXXXXXXXXXFW, S11 => XXDXXXXXXXXXXXXXXXFK, Y
                           => XXDXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXXWDXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXXXXXP, D1 => 
                           wp(1), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXQ, D3 => 
                           XXDXXXXXX, S00 => XXYPXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S11 => XXDXXXXXX, Y 
                           => axwdata(1));
   XXDXXXXXXXXXXXXWDXXXXXXXK : DFE3C port map( D => XXDXXXXXXXXXXHV, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXXXXXXXFF : OR2B port map( A => XXDDXXXXXP, B => 
                           XXDDXXXXXH, Y => XXDXXXXXXXXXXXXXXXXXXXXXXXXKP);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXJ : AND4A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFJ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFH);
   XXDXXXXXXXXXXXXXWXDDXXXXXP : CM8 port map( D0 => waddr(3), D1 => XXDDXXXXXP,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(3));
   XXDXXXXXXXXXXXXXXWXXXXXXXXXX : CM8INV port map( A => waddr(10), Y => 
                           XXDXXXXXXXXXXXXXXXWXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXL : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXF);
   XXDXXXXXXXXXXXXXXDDXXXXXK : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXK, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXW);
   XXDXXXXXXXXXXXXXXXDDXXXXXK : CM8 port map( D0 => raddr(9), D1 => XXDDXXXXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(9));
   XXDXXXXXXXXXXXXXWDXXXXXXXXFH : CM8 port map( D0 => wdata(6), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFQ, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(13));
   XXDXXXXXXXXXXXXXXXXXXXLXXFP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHJ, D1 => tmout(14),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D3 => 
                           tmout(14), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKD, S11 => XXDXXXXXX, Y 
                           => XXDXXXXXXXXXXXXXXXXXXXXLXXXHF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXJ : CM8 port map( D0 => XXDXXXXXXXXXXJK, D1 => 
                           axrdata(13), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(6));
   XXDXXXXXXXXXXXXXWDXXXXXXXXFJ : CM8 port map( D0 => wdata(13), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFK, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(20));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, S01 => VXXXXXXXX,
                           S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD);
   XXDXXXXXXXXXXXXXXXXXXXLXXFQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHL, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D2 => tmout(33), D3 
                           => tmout(33), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHL, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S10 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S11 => XXDXXXXXX, 
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S01 => VXXXXXXXX,
                           S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXL, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFW);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFL : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXV);
   XXDXXXXXXXXXXXXXXDDX : DFE3C port map( D => XXDXXXXXXXXXXXXXXXXX, E => 
                           XXDXXXXXXXXXXYXXL, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXDDXX);
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXX : OR3A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, B => 
                           XXDXXXXXXXXXXXXXXXXXF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX);
   XXDXXXXXXXXXXXXXWXDDXXXXXQ : CM8 port map( D0 => waddr(2), D1 => XXDDXXXXXQ,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(2));
   XXDXXXXXXXXXXXXXWDXXXXXXXXFK : CM8 port map( D0 => wdata(5), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXJ, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(12));
   XXDXXXXXXXXXXXXXWDXXXXXXXXFL : CM8 port map( D0 => wdata(14), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXK, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(21));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHK);
   XXDXXXXXXXXXXXXXXXXXXXLXXFV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHP, D1 => tmout(28),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, D3 => 
                           tmout(28), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJD);
   XXDXXXXXXXXXXXXXXXK : XOR2 port map( A => XXDDXXXXXL, B => waddr(4), Y => 
                           XXDXXXXXXXXXXXXXXXFW);
   XXDXXXXXXXXXXXXXXXDDXXXXXL : CM8 port map( D0 => raddr(8), D1 => XXDDXXXXXF,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(8));
   XXDXXXXXXXXXXXXXXDDXXXXXL : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXP, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXV);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXF, D1 => 
                           axrdata(14), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(7));
   XXDXXXXXXXXXXXXXWDXXXXXXXL : CM8 port map( D0 => XXDXXXXXXXXXXXXXXL, D1 => 
                           wp(0), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXX, D3 => 
                           XXDXXXXXX, S00 => XXYPXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S11 => XXDXXXXXX, Y 
                           => axwdata(0));
   XXDXXXXXXXXXXXXWDXXXXXXXL : DFE3C port map( D => XXDXXXXXXXXXXFV, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXF,
                           D1 => VXXXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX
                           );
   XXDXXXXXXXXXXXXWDXXXXXXXXFK : DFE3C port map( D => XXDXXXXXXXXXXHQ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHF);
   XXDXXXXXXXXXXXXWDXXXXXXXXFL : DFE3C port map( D => XXDXXXXXXXXXXP, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXX, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHH : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXK, E => XXDXXXXXXXXXXYXXK
                           , CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXYXXJ, D2 => XXDXXXXXX, D3 => XXDXXXXXX,
                           S00 => XXDXXXXXXXXXXYXX, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXW, S11 => XXDXXXXXXXXXXXXXXXHJ, Y 
                           => XXDXXXXXXXXXXYXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXXXXXXXXXXXXXDX, D2 => VXXXXXXXX, D3 => VXXXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, S10 => 
                           XXDXXXXXXXXXXXXXXXFJ, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXXXXFLXXXXXXX : AND3A port map( A => XXXXXXDXXXX, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXFLXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHW, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJJ);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXJ, D1 => VXXXXXXXX, D2 => 
                           XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXF, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXX, S11 => 
                           XXDXXXXXXXXXXY, Y => XXDXXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXV, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJD, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           VXXXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXXXXXXY, 
                           S00 => XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX, S01 =>
                           XXDXXXXXXXXXXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXJ, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXYXXF);
   XXDXXXXXXXXXXXXWDXXXXXXXP : DFE3C port map( D => XXDXXXXXXXXXXHF, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFK);
   XXDXXXXXXXXXXXXXXXL : XOR2 port map( A => XXDDXXXXXF, B => rds(0), Y => 
                           XXDXXXXXXXXXXXXXXXHV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXQ, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFV : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHP);
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXXXXXXYXXQ,
                           D1 => XXDXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, 
                           S00 => XXDXXXXXXXXXXXXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, S11 => 
                           XXDXXXXXXXXXXYXXV, Y => XXDXXXXXXXXXXYXXL);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D2 => VXXXXXXXX, 
                           D3 => VXXXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXX, S01 
                           => XXDXXXXXXXXXXXXXXXFH, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, S11 => XXDXXXXXX, 
                           Y => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXX, D1 => tmout(5), D2 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, D3 => tmout(5)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH
                           , S11 => XXDXXXXXXXXXXXXXXXXXXXXXXXFJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXFW : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFV);
   XXDXXXXXXXXXXXXXDDXXLXP : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXH, S00 => XXDDXXXXXK, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXF, 
                           S11 => XXDXXXXXXXXXXYXXXK, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXFW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFW, D1 => tmout(21),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, D3 => 
                           tmout(21), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKF, S11 => XXDXXXXXX, Y 
                           => XXDXXXXXXXXXXXXXXXXXXXXLXXXHV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHL : AND3B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXWDXXXXXXXXFP : DFE3C port map( D => XXDXXXXXXXXXXFP, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXWDXXXXXXXXFQ : DFE3C port map( D => XXDXXXXXXXXXXHJ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHD : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXJ);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXX : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXF, D1 => VXXXXXXXX, D2 => 
                           XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX);
   XXDXXXXXXXXXXXXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXXHQ, E => 
                           XXDXXXXXXXXXXYXXH, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXFH);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXX : AND2A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXF, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXDDXXLXX : XA1 port map( A => XXDXXXXXXXXXXXXXXDDXXXXXFJ, B 
                           => XXDDXXXXXXF, C => XXDXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXDXXXXX : AND2 port map( A => XXDXXXXXXXXXXXXWXX, 
                           B => XXDXXXXXXXXXXXXXXDDXXXXXFD, Y => 
                           XXXXXXXXXXXXXXDX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHJ, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHK, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXX : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXLXQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXJ, D1 => tmout(2), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, D3 => 
                           tmout(2), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 
                           => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXFD, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXK);
   XXDXXXXXXXXXXXXXDDXLDXXX : CM8 port map( D0 => VXXXXXXXX, D1 => XXDXXXXXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXLDXXXXXXXXX, S01 => 
                           XXDXXXXXXXXXXYXXJ, S10 => XXDXXXXXXXXXXYXXV, S11 => 
                           XXDXXXXXXXXXXYXXW, Y => XXDXXXXXXXXXXXXXDDXXF);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXX : OR2 port map( A => 
                           XXDXXXXXXXXXXXFXXXXLXXDX, B => stop_scrub, Y => 
                           XXDXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXPXXXXJ : CM8 port map( D0 => XXDXXXXXXXXXXJV, D1 => 
                           axrdata(4), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rp(4));
   XXDXXXXXXXXXXXXXXXXXXXLXXHD : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHF, D1 => tmout(26),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHK, D3 => 
                           tmout(26), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXFF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXPXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXHF, D1 => 
                           axrdata(5), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rp(5));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXL : CM8INV port map( A => axrdata(10), Y => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXDDXXLXQ : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXH, S00 => XXDXXXXXXXXXXXXXXXFP, 
                           S01 => VXXXXXXXX, S10 => XXDDXXXXXQ, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXDDXXLXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXP);
   XXDXXXXXXXXXXXXXDDXXXXXF : NAND4 port map( A => XXDDXXXXXW, B => XXDDXXXXXV,
                           C => XXDDXXXXXQ, D => XXDDXXXXXP, Y => 
                           XXDXXXXXXXXXXYXXXK);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXLXXHF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFV, D1 => tmout(13),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, D3 => 
                           tmout(13), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXH, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXQ, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH);
   XXDXXXXXXXXXXXXXXXXXXLDXXXXXXXX : AND4B port map( A => XXXXXXDXXXX, B => 
                           XXDXXXXXXXXXXXXXXXXXF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXWXXXXXX : CM8 port map( D0 => we, D1 => XXDXXXXXXXXXXXXWXX, 
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFD, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwe);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXV : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXH);
   XXDXXXXXXXXXXXXXDDXXXXL : AND2A port map( A => XXYPXXXXXXF, B => 
                           XXDXXXXXXXXXXXXXXXHK, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXHW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXP, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ : AND3B port map( A => XXXXXXXXXLXXF, B 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXHJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXFH : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, D2 => VXXXXXXXX
                           , D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKV);
   XXDXXXXXXXXXXXXXXXXXXXXXXFJ : OR3 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKW, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJH, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXFK : OR4 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLH, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKQ);
   XXDXXXXXXXXXXXXXXXXXXXLXXHH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHQ, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, D2 => tmout(41)
                           , D3 => tmout(41), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLF, S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXXFP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFL, D1 => XXDXXXXXX, 
                           D2 => wdata(28), D3 => XXDXXXXXX, S00 => XXDXXXXXX, 
                           S01 => XXDXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXWDXXXXXXXXXXXXXXXXXXX, S11 => 
                           XXYPXXXXXX, Y => axwdata(35));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXW : CM8 port map( D0 => XXDXXXXXXXXXXL, D1 => 
                           axrdata(30), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXF, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(23));
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           waddr(7), Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXWDXXXXXXXQ : DFE3C port map( D => XXDXXXXXXXXXXJV, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFD : CM8 port map( D0 => axrdata(17), D1 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXJ, D2 => 
                           axrdata(17), D3 => axrdata(17), S00 => 
                           XXDXXXXXXXXXXV, S01 => XXDXXXXXXXXXXH, S10 => 
                           XXYPXXXXXXH, S11 => XXDXXXXXXXXF, Y => rdata(10));
   XXDXXXXXXXXXXXXXXXDDXXXXXP : CM8 port map( D0 => raddr(5), D1 => XXDDXXXXXK,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(5));
   XXDXXXXXXXXXXXXXXXXXXXLXXHJ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXJ, D1 => tmout(34), D2 
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXLH, D3 => tmout(34), 
                           S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S01 => 
                           VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXV);
   XXDXXXXXXXXXXXXXXXDDXXXXXQ : CM8 port map( D0 => raddr(4), D1 => XXDDXXXXXL,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(4));
   XXDXXXXXXXXXXXXXXXXXXXXXK : OR3 port map( A => XXDXXXXXXXXXXXXXXXXXXXXXXXFJ,
                           B => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXP, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXF : OR3A port map( A => 
                           XXDXXXXXXXXXXXXXXXDDXX, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLK, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLV, Y => 
                           XXDXXXXXXXXXXYXXQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXFL : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXFP, D2 => VXXXXXXXX, D3 => 
                           VXXXXXXXX, S00 => XXDDXXXXXK, S01 => XXDDXXXXXJ, S10
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXKP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLV);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFF : CM8 port map( D0 => XXDXXXXXXXXXXJQ, D1 =>
                           axrdata(18), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(11));
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHK : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXK);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFH : CM8 port map( D0 => axrdata(29), D1 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXX, D2 => 
                           axrdata(29), D3 => axrdata(29), S00 => 
                           XXDXXXXXXXXXXV, S01 => XXDXXXXXXXXXXJF, S10 => 
                           XXYPXXXXXXF, S11 => XXDXXXXXXXX, Y => rdata(22));
   XXDXXXXXXXXXXXXXDDXXXXP : AND2A port map( A => XXYPXXXXXXF, B => 
                           XXDXXXXXXXXXXXXXXXHK, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH);
   XXDXXXXXXXXXXXXWDXXXXXXXXFV : DFE3C port map( D => XXDXXXXXXXXXXHD, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXW);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXJ : CM8INV port map( A => axrdata(35), Y 
                           => XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHL : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHP : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHD);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFL);
   XXDXXXXXXXXXXXXXWDXXXXXXXXFQ : CM8 port map( D0 => wdata(27), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXP, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(34));
   XXDXXXXXXXXXXXXWDXXXXXXXXFW : DFE3C port map( D => XXDXXXXXXXXXXF, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFH);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX : OR2 port map( A => 
                           XXDXXXXXXXXXXXFXXXXLXXDX, B => stop_scrub, Y => 
                           XXDXXXXXXXXXXYXXV);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : AND4A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, B => 
                           XXDXXXXXXXXXXXXXXXFH, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, D => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXHL);
   XXDXXXXXXXXXXXXXXXXXXXXXXFP : OR4B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXL, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXJ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLP);
   XXDXXXXXXXXXXXXXDDXXLXV : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXH, S00 => XXDDXXXXXP, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXDDXXLXXXXXXXH, 
                           S11 => XXDXXXXXXXXXXXXXXXFP, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXW);
   XXDXXXXXXXXXXXXDXXXXXXXJ : CM8 port map( D0 => axrdata(10), D1 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXK, D2 => 
                           axrdata(10), D3 => axrdata(10), S00 => 
                           XXDXXXXXXXXXXV, S01 => XXDXXXXXXXXXXH, S10 => 
                           XXYPXXXXXX, S11 => XXDXXXXXXXX, Y => rdata(3));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJD : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHL, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV);
   XXDXXXXXXXXXXXXXXDDXXXXXX : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXXF,
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXX);
   XXDXXXXXXXXXXXXDXXXXXXXK : CM8 port map( D0 => XXDXXXXXXXXXXFV, D1 => 
                           axrdata(9), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXYPXXXXXX, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 
                           => XXDXXXXXX, Y => rdata(2));
   XXDXXXXXXXXXXXXXXDDXXXXXXF : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXX,
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXXF);
   XXDXXXXXXXXXXXXXXXP : XOR2 port map( A => XXDDXXXXX, B => rds(1), Y => 
                           XXDXXXXXXXXXXXXXXXFL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJF : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXV, E => XXDXXXXXXXXXXYXXK
                           , CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV);
   XXDXXXXXXXXXXXXXXXXXXXLXXHK : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHH, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D2 => tmout(27),
                           D3 => tmout(27), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKK, S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXHH);
   XXDXXXXXXXXXXXXXWXDDXXXXXV : CM8 port map( D0 => waddr(6), D1 => XXDDXXXXXJ,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(6));
   XXDXXXXXXXXXXXXXXXXXXLDXXXXXX : AND4B port map( A => XXXXXXDXXXX, B => 
                           XXDXXXXXXXXXXYXXV, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXYXXK);
   XXDXXXXXXXXXXXXXXXXXXXLXV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXH, D1 => tmout(3), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, D3 => tmout(3)
                           , S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV
                           , S11 => XXDXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXL);
   XXDXXXXXXXXXXXXWDXXXXXXXXHD : DFE3C port map( D => XXDXXXXXXXXXXFK, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHD);
   XXDXXXXXXXXXXXXWDXXXXXXXXHF : DFE3C port map( D => XXDXXXXXXXXXXFJ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHK);
   XXDXXXXXXXXXXXXXXXXXXXLXXHL : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHK, D1 => tmout(15),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHH, D3 => 
                           tmout(15), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXW);
   XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXXXXXXF : OR3A port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, B => 
                           XXDXXXXXXXXXXXXXXXXXF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXWDXXXXXXXP : CM8 port map( D0 => XXDXXXXXXXXXXXXXXK, D1 => 
                           wp(4), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXF, D3 => 
                           XXDXXXXXX, S00 => XXYPXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S11 => XXDXXXXXX, Y 
                           => axwdata(4));
   XXDXXXXXXXXXXXXXXDDXXXXXP : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXQ, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFJ : CM8 port map( D0 => XXDXXXXXXXXXXFJ, D1 =>
                           axrdata(26), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(19));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXV : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD, D2 => VXXXXXXXX
                           , D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHP, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXXXXXXXLXXHP : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFL, D1 => tmout(12),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, D3 => 
                           tmout(12), S00 => XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX,
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKV, S11 => XXDXXXXXX, Y 
                           => XXDXXXXXXXXXXXXXXXXXXXXLXXXHQ);
   XXDXXXXXXXXXXXXXWDXXXXXXXXFV : CM8 port map( D0 => wdata(18), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXH, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(25));
   XXDXXXXXXXXXXXXXWXDDXXXXXX : CM8 port map( D0 => waddr(10), D1 => 
                           XXDDXXXXXXF, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S01 => VXXXXXXXX, S10
                           => XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(10));
   XXDXXXXXXXXXXXXXXXXXXLDXXXXXXXXF : AND4B port map( A => XXXXXXDXXXX, B => 
                           XXDXXXXXXXXXXXXXXXXXF, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, Y => 
                           XXDXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXXWDXXXXXXXXFW : CM8 port map( D0 => wdata(9), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXL, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(16));
   XXDXXXXXXXXXXXXXXXXXXXLXXHQ : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFQ, D1 => tmout(35),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHV, D3 => 
                           tmout(35), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKH, S11 => XXDXXXXXX, Y 
                           => XXDXXXXXXXXXXXXXXXXXXXXLXXXHL);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXX : CM8INV port map( A => XXXXXXDXXXX,
                           Y => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXWDXXXXXXXXHD : CM8 port map( D0 => wdata(17), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFV, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(24));
   XXDXXXXXXXXXXXXXDDXXXXXXXXXF : CM8INV port map( A => XXDXXXXXXXXXXYXXXK, Y 
                           => XXDXXXXXXXXXXXXXXDDXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, D2 => VXXXXXXXX
                           , D3 => VXXXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXF, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHQ, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFQ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXWDXXXXXXXXHF : CM8 port map( D0 => wdata(10), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFJ, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFL, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(17));
   XXDXXXXXXXXXXXXXXXQ : XOR2 port map( A => XXDDXXXXXQ, B => waddr(2), Y => 
                           XXDXXXXXXXXXXXXXXXHH);
   XXDXXXXXXXXXXXXXWDXXXXXXXXHH : CM8 port map( D0 => wdata(23), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXF, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(30));
   XXDXXXXXXXXXXXXXWDXXXXXXXQ : CM8 port map( D0 => XXDXXXXXXXXXXXXXXJ, D1 => 
                           wp(5), D2 => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXP, D3 => 
                           XXDXXXXXX, S00 => XXYPXXXXXX, S01 => VXXXXXXXX, S10 
                           => XXDXXXXXXXXXXXXXXDDXXXXXFF, S11 => XXDXXXXXX, Y 
                           => axwdata(5));
   XXDXXXXXXXXXXXXXXXXXXXLXXHV : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLD, D1 => tmout(40), D2 
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJF);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFK : CM8 port map( D0 => XXDXXXXXXXXXXJD, D1 =>
                           axrdata(25), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(18));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH);
   XXDXXXXXXXXXXXXXWXDDXXXXXW : CM8 port map( D0 => waddr(7), D1 => XXDDXXXXXH,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFH, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(7));
   XXDXXXXXXXXXXXXXWXDDXXXXXXF : CM8 port map( D0 => waddr(11), D1 => 
                           XXDDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           XXDXXXXXXXXXXXXXXDDXXXXXFF, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axwaddr(11));
   XXDXXXXXXXXXXXXXXXXXXXXXXFQ : OR3 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKF, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHJ, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXKW);
   XXDXXXXXXXXXXXXXXDDXXXXXQ : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXH, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXL);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => we, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => VXXXXXXXX, S00 => 
                           we, S01 => XXDDXXXXXP, S10 => waddr(3), S11 => 
                           XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXWDXXXXXXXXHJ : CM8 port map( D0 => wdata(22), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFW, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(29));
   XXDXXXXXXXXXXXXXDDXXLXXXXXXF : CM8INV port map( A => XXDDXXXXXL, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXH : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLK, D1 => XXDXXXXXX, D2 
                           => VXXXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, S01 => VXXXXXXXX, 
                           S10 => XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXXX, 
                           S11 => XXDXXXXXXXXXXXXXXXXXXXXXXXXLV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXDDXXXXXV : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXJ, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXX);
   XXDXXXXXXXXXXXXXXXXFLXX : DFC1B port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => tmoutflg);
   XXDXXXXXXXXXXXXXXXXXXXLXXHW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHD, D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJK, D2 => tmout(29)
                           , D3 => tmout(29), S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLW, S01 => VXXXXXXXX, S10
                           => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXL);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFL : CM8 port map( D0 => axrdata(22), D1 => 
                           XXDXXXXXXXXXXXXDXXXXXXXXXXXXXXXXXXXXXXXXF, D2 => 
                           axrdata(22), D3 => axrdata(22), S00 => 
                           XXDXXXXXXXXXXV, S01 => XXDXXXXXXXXXXFD, S10 => 
                           XXYPXXXXXXH, S11 => XXDXXXXXXXXJ, Y => rdata(15));
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFP : CM8 port map( D0 => XXDXXXXXXXXXXFH, D1 =>
                           axrdata(33), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXF, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(26));
   XXDXXXXXXXXXXXXXXXV : XOR2 port map( A => XXDDXXXXXK, B => waddr(5), Y => 
                           XXDXXXXXXXXXXXXXXXFD);
   XXDXXXXXXXXXXXXXWDXXXXXXXV : CM8 port map( D0 => wdata(1), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXL, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(8));
   XXDXXXXXXXXXXXXXXXDDXXXXXV : CM8 port map( D0 => raddr(0), D1 => XXDDXXXXXW,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(0));
   XXDXXXXXXXXXXXXWDXXXXXXXV : DFE3C port map( D => XXDXXXXXXXXXXQ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJH : AND2B port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXV, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXHF, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXXXXLXW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXF, D1 => tmout(4), D2
                           => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFH, D3 => 
                           tmout(4), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXX, S01 
                           => VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXXXXXXXXXFJ, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXLXXH);
   XXDXXXXXXXXXXXXXXXXXXXXXXFV : OR2B port map( A => XXDDXXXXXQ, B => 
                           XXDDXXXXXL, Y => XXDXXXXXXXXXXXXXXXXXXXXXXXXLL);
   XXDXXXXXXXXXXXXXWDXXXXXXXW : CM8 port map( D0 => wdata(2), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXH, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFF, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(9));
   XXDXXXXXXXXXXXXWDXXXXXXXW : DFE3C port map( D => XXDXXXXXXXXXXJP, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXLXXJD : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, D1 => tmout(32),
                           D2 => XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXFP, D3 => 
                           tmout(32), S00 => XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF, 
                           S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S11 => XXDXXXXXX, 
                           Y => XXDXXXXXXXXXXXXXXXXXXXXLXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXXXL : OR4 port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ, B => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXW, C => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL, D => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFV, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFQ : CM8 port map( D0 => XXDXXXXXXXXXXJH, D1 =>
                           axrdata(34), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXF, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(27));
   XXDXXXXXXXXXXXXXXDDXXXXXW : DFE3C port map( D => XXDXXXXXXXXXXXXXXDDXXLXXL, 
                           E => XXDXXXXXXXXXXXXXDDXXF, CLK => clk, CLR => rstn,
                           Q => XXDDXXXXXF);
   XXDXXXXXXXXXXXXXXXDDXXXXXW : CM8 port map( D0 => raddr(1), D1 => XXDDXXXXXV,
                           D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXX, S01 => VXXXXXXXX, S10 => 
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axraddr(1));
   XXDXXXXXXXXXXXXXXXXXXXXXXFW : CM8 port map( D0 => XXDXXXXXX, D1 => VXXXXXXXX
                           , D2 => VXXXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXQ, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXH, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK, S11 => XXDXXXXXX
                           , Y => XXDXXXXXXXXXXXXXXXXXXXXXXXXKL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXW : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF, S01 => 
                           VXXXXXXXX, S10 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXK);
   XXDXXXXXXXXXXXXDXXXXXXXXXXXXXFV : CM8 port map( D0 => XXDXXXXXXXXXXFW, D1 =>
                           axrdata(21), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 
                           => XXYPXXXXXXH, S01 => VXXXXXXXX, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => rdata(14));
   XXDXXXXXXXXXXXXXWDXXXXXXXXHK : CM8 port map( D0 => wdata(21), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXX, D2 => XXDXXXXXX, D3
                           => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, S01
                           => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y 
                           => axwdata(28));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJJ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXH, E => XXDXXXXXXXXXXYXXK
                           , CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFF);
   XXDXXXXXXXXXXXXXWDXXXXXXXXHL : CM8 port map( D0 => wdata(24), D1 => 
                           XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXFP, D2 => XXDXXXXXX, 
                           D3 => XXDXXXXXX, S00 => XXDXXXXXXXXXXXXXXDDXXXXXFD, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => axwdata(31));
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJK : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJ, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJD);
   XXDXXXXXXXXXXXXXDDXXLXXF : CM8 port map( D0 => XXDXXXXXX, D1 => 
                           XXDXXXXXXXXXXXXXXXXXH, D2 => XXDXXXXXXXXXXXXXXXXXH, 
                           D3 => XXDXXXXXX, S00 => XXDDXXXXXXF, S01 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFJ, S10 => XXDDXXXXXX, S11 
                           => XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXDDXXLXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJL : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHP, E => 
                           XXDXXXXXXXXXXYXXK, CLK => clk, CLR => rstn, Q => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJP);
   XXDXXXXXXXXXXXXWDXXXXXXXXHH : DFE3C port map( D => XXDXXXXXXXXXXJQ, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHL);
   XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXF, D1 => VXXXXXXXX, D2 => 
                           XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXPXXXXXXXXXXF);
   XXDXXXXXXXXXXXXXXXXXXXXQXXXXXXXXF : CM8 port map( D0 => VXXXXXXXX, D1 => 
                           XXDXXXXXX, D2 => VXXXXXXXX, D3 => XXDXXXXXXXXXXXXWXX
                           , S00 => XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXDDXXX, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXXXXXXXXQXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXXXXXV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXF, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFJ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJP : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXF, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXJF);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXF : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFD, Y => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXX);
   XXDXXXXXXXXXXXXXXXXXXXH : CM8 port map( D0 => re, D1 => XXDXXXXXXXXXXXXXXXFH
                           , D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXDDXXXXXFD, S01 => VXXXXXXXX, S10 =>
                           XXDXXXXXX, S11 => XXDXXXXXX, Y => axre);
   XXDXXXXXXXXXXXXWDXXXXXXXXHJ : DFE3C port map( D => XXDXXXXXXXXXXFH, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXHH);
   XXDXXXXXXXXXXXXWDXXXXXXXXHK : DFE3C port map( D => XXDXXXXXXXXXXHP, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXXXXF, CLK => clk, CLR =>
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXV);
   XXDXXXXXXXXXXXXXDDXXLXXXXXXH : CM8INV port map( A => XXDDXXXXXQ, Y => 
                           XXDXXXXXXXXXXXXXXDDXXLXXXXXXXH);
   XXDXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXQXXXXXXXXXXXXXXXXXXXF, D1 => 
                           VXXXXXXXX, D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXK, S01 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXFF, S10 => XXDXXXXXX, 
                           S11 => XXDXXXXXX, Y => XXDXXXXXXXXXXYXXJ);
   XXDXXXXXXXXXXXXXDDXXLXW : CM8 port map( D0 => XXDXXXXXXXXXXXXXXXXXH, D1 => 
                           XXDXXXXXX, D2 => XXDXXXXXX, D3 => 
                           XXDXXXXXXXXXXXXXXXXXH, S00 => XXDXXXXXXXXXXYXXXK, 
                           S01 => VXXXXXXXX, S10 => XXDDXXXXXL, S11 => 
                           XXDXXXXXX, Y => XXDXXXXXXXXXXXXXXDDXXLXXH);
   XXDXXXXXXXXXXXXPXXXXL : CM8 port map( D0 => XXDXXXXXXXXXXJP, D1 => 
                           axrdata(0), D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 =>
                           bypass, S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => 
                           XXDXXXXXX, Y => rp(0));
   XXDXXXXXXXXXXXXXXXXXXXLXXJF : CM8 port map( D0 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLQ, D1 => tmout(20), D2 
                           => XXDXXXXXX, D3 => XXDXXXXXX, S00 => 
                           XXDXXXXXXXXXXXXXXXXXXPXXXXXXXXXXX, S01 => VXXXXXXXX,
                           S10 => XXDXXXXXX, S11 => XXDXXXXXX, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXJ);
   XXDXXXXXXXXXXXXPXXXXP : CM8 port map( D0 => XXDXXXXXXXXXXQ, D1 => axrdata(1)
                           , D2 => XXDXXXXXX, D3 => XXDXXXXXX, S00 => bypass, 
                           S01 => VXXXXXXXX, S10 => XXDXXXXXX, S11 => XXDXXXXXX
                           , Y => rp(1));
   XXDXXXXXXXXXXXXWDXXXXXXXXHL : DFE3C port map( D => XXDXXXXXXXXXX, E => 
                           XXDXXXXXXXXXXXXXXDDXXXXXQXXXX, CLK => clk, CLR => 
                           rstn, Q => XXDXXXXXXXXXXXXWDXXXXXXXXXXXXXXQ);
   XXDXXXXXXXXXXXXXXXXXXXXXXXW : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXW, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXL);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJQ : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHQ, E => 
                           XXDXXXXXXXXXXXXXXXXXK, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFP);
   XXDXXXXXXXXXXXXXXXXXXXXXXHD : CM8 port map( D0 => rds(2), D1 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXH, D2 => VXXXXXXXX, 
                           D3 => VXXXXXXXX, S00 => XXDDXXXXXXF, S01 => 
                           VXXXXXXXX, S10 => XXDXXXXXXXXXXXXXXXHV, S11 => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLJ, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXLK);
   XXDXXXXXXXXXXXXXXXXXXXXXXXXJV : DFE3C port map( D => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXHV, E => 
                           XXDXXXXXXXXXXXXXXXXXL, CLK => clk, CLR => rstn, Q =>
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFW);
   XXDXXXXXXXXXXXXXXXXXXXXXP : DFC1B port map( D => XXDXXXXXXXXXXYXXXJ, CLK => 
                           clk, CLR => rstn, Q => XXDXXXXXXXXXXXXXXXXXXXXXXXFH)
                           ;
   XXDXXXXXXXXXXXXXXXXXXXLXXXXXXXHQ : CM8INV port map( A => 
                           XXDXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXFK, Y => 
                           XXDXXXXXXXXXXXXXXXXXXXXLXXXXXXXXHQ);

end SYN_DEF_ARCH;
