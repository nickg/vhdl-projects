library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

--
entity oskmem is
  port (Clk : in std_logic;
        address : in integer range 0 to 4095;
        we : in std_logic;
        data_i : in unsigned(7 downto 0);
        data_o : out unsigned(7 downto 0);
        writes : out unsigned(7 downto 0);
        no_writes : out unsigned(7 downto 0)
        );
end oskmem;

architecture Behavioral of oskmem is

  signal write_count : unsigned(7 downto 0) := x"00";
  signal no_write_count : unsigned(7 downto 0) := x"00";
  
  type ram_t is array (0 to 4095) of unsigned(7 downto 0);
  constant initram : ram_t := (
          x"00", -- $00000
          x"00", -- $00001
          x"00", -- $00002
          x"00", -- $00003
          x"00", -- $00004
          x"00", -- $00005
          x"00", -- $00006
          x"00", -- $00007
          x"7c", -- $00008
          x"82", -- $00009
          x"aa", -- $0000a
          x"82", -- $0000b
          x"ba", -- $0000c
          x"82", -- $0000d
          x"7c", -- $0000e
          x"00", -- $0000f
          x"7c", -- $00010
          x"ba", -- $00011
          x"fe", -- $00012
          x"fe", -- $00013
          x"ba", -- $00014
          x"c6", -- $00015
          x"7c", -- $00016
          x"00", -- $00017
          x"6c", -- $00018
          x"fe", -- $00019
          x"fe", -- $0001a
          x"fe", -- $0001b
          x"7c", -- $0001c
          x"38", -- $0001d
          x"10", -- $0001e
          x"00", -- $0001f
          x"10", -- $00020
          x"38", -- $00021
          x"7c", -- $00022
          x"fe", -- $00023
          x"7c", -- $00024
          x"38", -- $00025
          x"10", -- $00026
          x"00", -- $00027
          x"10", -- $00028
          x"38", -- $00029
          x"54", -- $0002a
          x"ee", -- $0002b
          x"54", -- $0002c
          x"10", -- $0002d
          x"fe", -- $0002e
          x"00", -- $0002f
          x"10", -- $00030
          x"38", -- $00031
          x"7c", -- $00032
          x"fe", -- $00033
          x"fe", -- $00034
          x"38", -- $00035
          x"7c", -- $00036
          x"00", -- $00037
          x"00", -- $00038
          x"00", -- $00039
          x"10", -- $0003a
          x"38", -- $0003b
          x"10", -- $0003c
          x"00", -- $0003d
          x"00", -- $0003e
          x"00", -- $0003f
          x"00", -- $00040
          x"7c", -- $00041
          x"7c", -- $00042
          x"6c", -- $00043
          x"7c", -- $00044
          x"7c", -- $00045
          x"00", -- $00046
          x"00", -- $00047
          x"30", -- $00048
          x"48", -- $00049
          x"84", -- $0004a
          x"84", -- $0004b
          x"48", -- $0004c
          x"30", -- $0004d
          x"00", -- $0004e
          x"00", -- $0004f
          x"fe", -- $00050
          x"fe", -- $00051
          x"fe", -- $00052
          x"fe", -- $00053
          x"fe", -- $00054
          x"fe", -- $00055
          x"fe", -- $00056
          x"00", -- $00057
          x"00", -- $00058
          x"14", -- $00059
          x"08", -- $0005a
          x"34", -- $0005b
          x"f0", -- $0005c
          x"a0", -- $0005d
          x"e0", -- $0005e
          x"00", -- $0005f
          x"10", -- $00060
          x"28", -- $00061
          x"10", -- $00062
          x"38", -- $00063
          x"10", -- $00064
          x"10", -- $00065
          x"00", -- $00066
          x"00", -- $00067
          x"30", -- $00068
          x"38", -- $00069
          x"28", -- $0006a
          x"20", -- $0006b
          x"20", -- $0006c
          x"e0", -- $0006d
          x"c0", -- $0006e
          x"00", -- $0006f
          x"38", -- $00070
          x"48", -- $00071
          x"78", -- $00072
          x"48", -- $00073
          x"58", -- $00074
          x"d8", -- $00075
          x"c0", -- $00076
          x"00", -- $00077
          x"10", -- $00078
          x"5a", -- $00079
          x"24", -- $0007a
          x"66", -- $0007b
          x"24", -- $0007c
          x"5a", -- $0007d
          x"08", -- $0007e
          x"00", -- $0007f
          x"80", -- $00080
          x"e0", -- $00081
          x"f8", -- $00082
          x"fc", -- $00083
          x"f8", -- $00084
          x"e0", -- $00085
          x"80", -- $00086
          x"00", -- $00087
          x"04", -- $00088
          x"1c", -- $00089
          x"7c", -- $0008a
          x"fc", -- $0008b
          x"7c", -- $0008c
          x"1c", -- $0008d
          x"04", -- $0008e
          x"00", -- $0008f
          x"20", -- $00090
          x"70", -- $00091
          x"a8", -- $00092
          x"20", -- $00093
          x"a8", -- $00094
          x"70", -- $00095
          x"20", -- $00096
          x"00", -- $00097
          x"6c", -- $00098
          x"6c", -- $00099
          x"6c", -- $0009a
          x"6c", -- $0009b
          x"6c", -- $0009c
          x"00", -- $0009d
          x"6c", -- $0009e
          x"00", -- $0009f
          x"7c", -- $000a0
          x"e8", -- $000a1
          x"e8", -- $000a2
          x"68", -- $000a3
          x"28", -- $000a4
          x"28", -- $000a5
          x"28", -- $000a6
          x"00", -- $000a7
          x"1c", -- $000a8
          x"22", -- $000a9
          x"58", -- $000aa
          x"44", -- $000ab
          x"34", -- $000ac
          x"88", -- $000ad
          x"70", -- $000ae
          x"00", -- $000af
          x"00", -- $000b0
          x"00", -- $000b1
          x"fe", -- $000b2
          x"fe", -- $000b3
          x"00", -- $000b4
          x"00", -- $000b5
          x"00", -- $000b6
          x"00", -- $000b7
          x"10", -- $000b8
          x"38", -- $000b9
          x"54", -- $000ba
          x"10", -- $000bb
          x"54", -- $000bc
          x"38", -- $000bd
          x"7c", -- $000be
          x"00", -- $000bf
          x"30", -- $000c0
          x"78", -- $000c1
          x"fc", -- $000c2
          x"30", -- $000c3
          x"30", -- $000c4
          x"30", -- $000c5
          x"30", -- $000c6
          x"00", -- $000c7
          x"30", -- $000c8
          x"30", -- $000c9
          x"30", -- $000ca
          x"30", -- $000cb
          x"fc", -- $000cc
          x"78", -- $000cd
          x"30", -- $000ce
          x"00", -- $000cf
          x"08", -- $000d0
          x"0c", -- $000d1
          x"fe", -- $000d2
          x"fe", -- $000d3
          x"0c", -- $000d4
          x"08", -- $000d5
          x"00", -- $000d6
          x"00", -- $000d7
          x"20", -- $000d8
          x"60", -- $000d9
          x"fe", -- $000da
          x"fe", -- $000db
          x"60", -- $000dc
          x"20", -- $000dd
          x"00", -- $000de
          x"00", -- $000df
          x"c0", -- $000e0
          x"c0", -- $000e1
          x"c0", -- $000e2
          x"c0", -- $000e3
          x"c0", -- $000e4
          x"fe", -- $000e5
          x"fe", -- $000e6
          x"00", -- $000e7
          x"28", -- $000e8
          x"6c", -- $000e9
          x"fe", -- $000ea
          x"fe", -- $000eb
          x"6c", -- $000ec
          x"28", -- $000ed
          x"00", -- $000ee
          x"00", -- $000ef
          x"10", -- $000f0
          x"38", -- $000f1
          x"38", -- $000f2
          x"7c", -- $000f3
          x"7c", -- $000f4
          x"fe", -- $000f5
          x"fe", -- $000f6
          x"00", -- $000f7
          x"fe", -- $000f8
          x"7c", -- $000f9
          x"7c", -- $000fa
          x"38", -- $000fb
          x"38", -- $000fc
          x"10", -- $000fd
          x"10", -- $000fe
          x"00", -- $000ff
          x"00", -- $00100
          x"00", -- $00101
          x"00", -- $00102
          x"00", -- $00103
          x"00", -- $00104
          x"00", -- $00105
          x"00", -- $00106
          x"00", -- $00107
          x"30", -- $00108
          x"30", -- $00109
          x"30", -- $0010a
          x"30", -- $0010b
          x"30", -- $0010c
          x"00", -- $0010d
          x"30", -- $0010e
          x"00", -- $0010f
          x"66", -- $00110
          x"66", -- $00111
          x"66", -- $00112
          x"00", -- $00113
          x"00", -- $00114
          x"00", -- $00115
          x"00", -- $00116
          x"00", -- $00117
          x"6c", -- $00118
          x"6c", -- $00119
          x"fe", -- $0011a
          x"6c", -- $0011b
          x"fe", -- $0011c
          x"6c", -- $0011d
          x"6c", -- $0011e
          x"00", -- $0011f
          x"30", -- $00120
          x"7c", -- $00121
          x"c0", -- $00122
          x"78", -- $00123
          x"0c", -- $00124
          x"f8", -- $00125
          x"30", -- $00126
          x"00", -- $00127
          x"c4", -- $00128
          x"cc", -- $00129
          x"18", -- $0012a
          x"30", -- $0012b
          x"60", -- $0012c
          x"cc", -- $0012d
          x"8c", -- $0012e
          x"00", -- $0012f
          x"78", -- $00130
          x"cc", -- $00131
          x"78", -- $00132
          x"70", -- $00133
          x"ce", -- $00134
          x"cc", -- $00135
          x"7e", -- $00136
          x"00", -- $00137
          x"06", -- $00138
          x"0c", -- $00139
          x"18", -- $0013a
          x"00", -- $0013b
          x"00", -- $0013c
          x"00", -- $0013d
          x"00", -- $0013e
          x"00", -- $0013f
          x"18", -- $00140
          x"30", -- $00141
          x"60", -- $00142
          x"60", -- $00143
          x"60", -- $00144
          x"30", -- $00145
          x"18", -- $00146
          x"00", -- $00147
          x"60", -- $00148
          x"30", -- $00149
          x"18", -- $0014a
          x"18", -- $0014b
          x"18", -- $0014c
          x"30", -- $0014d
          x"60", -- $0014e
          x"00", -- $0014f
          x"00", -- $00150
          x"6c", -- $00151
          x"38", -- $00152
          x"fe", -- $00153
          x"38", -- $00154
          x"6c", -- $00155
          x"00", -- $00156
          x"00", -- $00157
          x"00", -- $00158
          x"30", -- $00159
          x"30", -- $0015a
          x"fc", -- $0015b
          x"30", -- $0015c
          x"30", -- $0015d
          x"00", -- $0015e
          x"00", -- $0015f
          x"00", -- $00160
          x"00", -- $00161
          x"00", -- $00162
          x"00", -- $00163
          x"30", -- $00164
          x"30", -- $00165
          x"60", -- $00166
          x"00", -- $00167
          x"00", -- $00168
          x"00", -- $00169
          x"00", -- $0016a
          x"7c", -- $0016b
          x"00", -- $0016c
          x"00", -- $0016d
          x"00", -- $0016e
          x"00", -- $0016f
          x"00", -- $00170
          x"00", -- $00171
          x"00", -- $00172
          x"00", -- $00173
          x"00", -- $00174
          x"30", -- $00175
          x"30", -- $00176
          x"00", -- $00177
          x"04", -- $00178
          x"0c", -- $00179
          x"18", -- $0017a
          x"30", -- $0017b
          x"60", -- $0017c
          x"c0", -- $0017d
          x"80", -- $0017e
          x"00", -- $0017f
          x"78", -- $00180
          x"cc", -- $00181
          x"dc", -- $00182
          x"fc", -- $00183
          x"ec", -- $00184
          x"cc", -- $00185
          x"78", -- $00186
          x"00", -- $00187
          x"30", -- $00188
          x"70", -- $00189
          x"30", -- $0018a
          x"30", -- $0018b
          x"30", -- $0018c
          x"30", -- $0018d
          x"fc", -- $0018e
          x"00", -- $0018f
          x"78", -- $00190
          x"cc", -- $00191
          x"0c", -- $00192
          x"38", -- $00193
          x"60", -- $00194
          x"c0", -- $00195
          x"fc", -- $00196
          x"00", -- $00197
          x"78", -- $00198
          x"cc", -- $00199
          x"0c", -- $0019a
          x"18", -- $0019b
          x"0c", -- $0019c
          x"cc", -- $0019d
          x"78", -- $0019e
          x"00", -- $0019f
          x"0c", -- $001a0
          x"1c", -- $001a1
          x"3c", -- $001a2
          x"cc", -- $001a3
          x"fe", -- $001a4
          x"0c", -- $001a5
          x"0c", -- $001a6
          x"00", -- $001a7
          x"fc", -- $001a8
          x"c0", -- $001a9
          x"f8", -- $001aa
          x"0c", -- $001ab
          x"0c", -- $001ac
          x"8c", -- $001ad
          x"78", -- $001ae
          x"00", -- $001af
          x"78", -- $001b0
          x"cc", -- $001b1
          x"c0", -- $001b2
          x"f8", -- $001b3
          x"cc", -- $001b4
          x"cc", -- $001b5
          x"78", -- $001b6
          x"00", -- $001b7
          x"fc", -- $001b8
          x"cc", -- $001b9
          x"18", -- $001ba
          x"30", -- $001bb
          x"30", -- $001bc
          x"30", -- $001bd
          x"30", -- $001be
          x"00", -- $001bf
          x"78", -- $001c0
          x"cc", -- $001c1
          x"cc", -- $001c2
          x"78", -- $001c3
          x"cc", -- $001c4
          x"cc", -- $001c5
          x"78", -- $001c6
          x"00", -- $001c7
          x"78", -- $001c8
          x"cc", -- $001c9
          x"cc", -- $001ca
          x"7c", -- $001cb
          x"0c", -- $001cc
          x"cc", -- $001cd
          x"78", -- $001ce
          x"00", -- $001cf
          x"00", -- $001d0
          x"30", -- $001d1
          x"30", -- $001d2
          x"00", -- $001d3
          x"30", -- $001d4
          x"30", -- $001d5
          x"00", -- $001d6
          x"00", -- $001d7
          x"00", -- $001d8
          x"30", -- $001d9
          x"30", -- $001da
          x"00", -- $001db
          x"30", -- $001dc
          x"30", -- $001dd
          x"60", -- $001de
          x"00", -- $001df
          x"00", -- $001e0
          x"18", -- $001e1
          x"30", -- $001e2
          x"60", -- $001e3
          x"30", -- $001e4
          x"18", -- $001e5
          x"00", -- $001e6
          x"00", -- $001e7
          x"00", -- $001e8
          x"00", -- $001e9
          x"7c", -- $001ea
          x"00", -- $001eb
          x"7c", -- $001ec
          x"00", -- $001ed
          x"00", -- $001ee
          x"00", -- $001ef
          x"00", -- $001f0
          x"30", -- $001f1
          x"18", -- $001f2
          x"0c", -- $001f3
          x"18", -- $001f4
          x"30", -- $001f5
          x"00", -- $001f6
          x"00", -- $001f7
          x"78", -- $001f8
          x"cc", -- $001f9
          x"0c", -- $001fa
          x"18", -- $001fb
          x"30", -- $001fc
          x"00", -- $001fd
          x"30", -- $001fe
          x"00", -- $001ff
          x"78", -- $00200
          x"cc", -- $00201
          x"dc", -- $00202
          x"dc", -- $00203
          x"c0", -- $00204
          x"cc", -- $00205
          x"78", -- $00206
          x"00", -- $00207
          x"30", -- $00208
          x"78", -- $00209
          x"cc", -- $0020a
          x"fc", -- $0020b
          x"cc", -- $0020c
          x"cc", -- $0020d
          x"cc", -- $0020e
          x"00", -- $0020f
          x"f8", -- $00210
          x"cc", -- $00211
          x"cc", -- $00212
          x"f8", -- $00213
          x"cc", -- $00214
          x"cc", -- $00215
          x"f8", -- $00216
          x"00", -- $00217
          x"78", -- $00218
          x"cc", -- $00219
          x"cc", -- $0021a
          x"c0", -- $0021b
          x"c0", -- $0021c
          x"cc", -- $0021d
          x"78", -- $0021e
          x"00", -- $0021f
          x"f0", -- $00220
          x"d8", -- $00221
          x"cc", -- $00222
          x"cc", -- $00223
          x"cc", -- $00224
          x"d8", -- $00225
          x"f0", -- $00226
          x"00", -- $00227
          x"fc", -- $00228
          x"c0", -- $00229
          x"c0", -- $0022a
          x"f0", -- $0022b
          x"c0", -- $0022c
          x"c0", -- $0022d
          x"fc", -- $0022e
          x"00", -- $0022f
          x"fc", -- $00230
          x"c0", -- $00231
          x"c0", -- $00232
          x"f0", -- $00233
          x"c0", -- $00234
          x"c0", -- $00235
          x"c0", -- $00236
          x"00", -- $00237
          x"78", -- $00238
          x"cc", -- $00239
          x"c0", -- $0023a
          x"dc", -- $0023b
          x"cc", -- $0023c
          x"cc", -- $0023d
          x"78", -- $0023e
          x"00", -- $0023f
          x"cc", -- $00240
          x"cc", -- $00241
          x"cc", -- $00242
          x"fc", -- $00243
          x"cc", -- $00244
          x"cc", -- $00245
          x"cc", -- $00246
          x"00", -- $00247
          x"fc", -- $00248
          x"30", -- $00249
          x"30", -- $0024a
          x"30", -- $0024b
          x"30", -- $0024c
          x"30", -- $0024d
          x"fc", -- $0024e
          x"00", -- $0024f
          x"3c", -- $00250
          x"18", -- $00251
          x"18", -- $00252
          x"18", -- $00253
          x"18", -- $00254
          x"d8", -- $00255
          x"70", -- $00256
          x"00", -- $00257
          x"cc", -- $00258
          x"d8", -- $00259
          x"f0", -- $0025a
          x"f0", -- $0025b
          x"f0", -- $0025c
          x"d8", -- $0025d
          x"cc", -- $0025e
          x"00", -- $0025f
          x"c0", -- $00260
          x"c0", -- $00261
          x"c0", -- $00262
          x"c0", -- $00263
          x"c0", -- $00264
          x"c0", -- $00265
          x"fc", -- $00266
          x"00", -- $00267
          x"c6", -- $00268
          x"ee", -- $00269
          x"fe", -- $0026a
          x"fe", -- $0026b
          x"d6", -- $0026c
          x"c6", -- $0026d
          x"c6", -- $0026e
          x"00", -- $0026f
          x"cc", -- $00270
          x"cc", -- $00271
          x"ec", -- $00272
          x"fc", -- $00273
          x"dc", -- $00274
          x"cc", -- $00275
          x"cc", -- $00276
          x"00", -- $00277
          x"78", -- $00278
          x"cc", -- $00279
          x"cc", -- $0027a
          x"cc", -- $0027b
          x"cc", -- $0027c
          x"cc", -- $0027d
          x"78", -- $0027e
          x"00", -- $0027f
          x"f8", -- $00280
          x"cc", -- $00281
          x"cc", -- $00282
          x"f8", -- $00283
          x"c0", -- $00284
          x"c0", -- $00285
          x"c0", -- $00286
          x"00", -- $00287
          x"78", -- $00288
          x"cc", -- $00289
          x"cc", -- $0028a
          x"cc", -- $0028b
          x"cc", -- $0028c
          x"78", -- $0028d
          x"0c", -- $0028e
          x"00", -- $0028f
          x"f8", -- $00290
          x"cc", -- $00291
          x"cc", -- $00292
          x"f8", -- $00293
          x"f0", -- $00294
          x"d8", -- $00295
          x"cc", -- $00296
          x"00", -- $00297
          x"78", -- $00298
          x"cc", -- $00299
          x"c0", -- $0029a
          x"78", -- $0029b
          x"0c", -- $0029c
          x"cc", -- $0029d
          x"78", -- $0029e
          x"00", -- $0029f
          x"fc", -- $002a0
          x"30", -- $002a1
          x"30", -- $002a2
          x"30", -- $002a3
          x"30", -- $002a4
          x"30", -- $002a5
          x"30", -- $002a6
          x"00", -- $002a7
          x"cc", -- $002a8
          x"cc", -- $002a9
          x"cc", -- $002aa
          x"cc", -- $002ab
          x"cc", -- $002ac
          x"cc", -- $002ad
          x"78", -- $002ae
          x"00", -- $002af
          x"cc", -- $002b0
          x"cc", -- $002b1
          x"cc", -- $002b2
          x"cc", -- $002b3
          x"cc", -- $002b4
          x"78", -- $002b5
          x"30", -- $002b6
          x"00", -- $002b7
          x"c6", -- $002b8
          x"c6", -- $002b9
          x"d6", -- $002ba
          x"fe", -- $002bb
          x"fe", -- $002bc
          x"ee", -- $002bd
          x"c6", -- $002be
          x"00", -- $002bf
          x"cc", -- $002c0
          x"cc", -- $002c1
          x"78", -- $002c2
          x"30", -- $002c3
          x"78", -- $002c4
          x"cc", -- $002c5
          x"cc", -- $002c6
          x"00", -- $002c7
          x"cc", -- $002c8
          x"cc", -- $002c9
          x"cc", -- $002ca
          x"78", -- $002cb
          x"30", -- $002cc
          x"30", -- $002cd
          x"30", -- $002ce
          x"00", -- $002cf
          x"fc", -- $002d0
          x"0c", -- $002d1
          x"18", -- $002d2
          x"30", -- $002d3
          x"60", -- $002d4
          x"e0", -- $002d5
          x"fc", -- $002d6
          x"00", -- $002d7
          x"78", -- $002d8
          x"60", -- $002d9
          x"60", -- $002da
          x"60", -- $002db
          x"60", -- $002dc
          x"60", -- $002dd
          x"78", -- $002de
          x"00", -- $002df
          x"00", -- $002e0
          x"80", -- $002e1
          x"c0", -- $002e2
          x"60", -- $002e3
          x"30", -- $002e4
          x"18", -- $002e5
          x"0c", -- $002e6
          x"00", -- $002e7
          x"78", -- $002e8
          x"18", -- $002e9
          x"18", -- $002ea
          x"18", -- $002eb
          x"18", -- $002ec
          x"18", -- $002ed
          x"78", -- $002ee
          x"00", -- $002ef
          x"10", -- $002f0
          x"38", -- $002f1
          x"6c", -- $002f2
          x"00", -- $002f3
          x"00", -- $002f4
          x"00", -- $002f5
          x"00", -- $002f6
          x"00", -- $002f7
          x"00", -- $002f8
          x"00", -- $002f9
          x"00", -- $002fa
          x"00", -- $002fb
          x"00", -- $002fc
          x"00", -- $002fd
          x"00", -- $002fe
          x"ff", -- $002ff
          x"c0", -- $00300
          x"60", -- $00301
          x"30", -- $00302
          x"00", -- $00303
          x"00", -- $00304
          x"00", -- $00305
          x"00", -- $00306
          x"00", -- $00307
          x"00", -- $00308
          x"00", -- $00309
          x"78", -- $0030a
          x"0c", -- $0030b
          x"7c", -- $0030c
          x"cc", -- $0030d
          x"7c", -- $0030e
          x"00", -- $0030f
          x"00", -- $00310
          x"60", -- $00311
          x"60", -- $00312
          x"7c", -- $00313
          x"66", -- $00314
          x"66", -- $00315
          x"7c", -- $00316
          x"00", -- $00317
          x"00", -- $00318
          x"00", -- $00319
          x"3c", -- $0031a
          x"60", -- $0031b
          x"60", -- $0031c
          x"60", -- $0031d
          x"3c", -- $0031e
          x"00", -- $0031f
          x"00", -- $00320
          x"06", -- $00321
          x"06", -- $00322
          x"3e", -- $00323
          x"66", -- $00324
          x"66", -- $00325
          x"3e", -- $00326
          x"00", -- $00327
          x"00", -- $00328
          x"00", -- $00329
          x"3c", -- $0032a
          x"66", -- $0032b
          x"7e", -- $0032c
          x"60", -- $0032d
          x"3c", -- $0032e
          x"00", -- $0032f
          x"00", -- $00330
          x"0e", -- $00331
          x"18", -- $00332
          x"3e", -- $00333
          x"18", -- $00334
          x"18", -- $00335
          x"18", -- $00336
          x"00", -- $00337
          x"00", -- $00338
          x"00", -- $00339
          x"3e", -- $0033a
          x"66", -- $0033b
          x"66", -- $0033c
          x"3e", -- $0033d
          x"06", -- $0033e
          x"7c", -- $0033f
          x"00", -- $00340
          x"60", -- $00341
          x"60", -- $00342
          x"7c", -- $00343
          x"66", -- $00344
          x"66", -- $00345
          x"66", -- $00346
          x"00", -- $00347
          x"00", -- $00348
          x"18", -- $00349
          x"00", -- $0034a
          x"38", -- $0034b
          x"18", -- $0034c
          x"18", -- $0034d
          x"3c", -- $0034e
          x"00", -- $0034f
          x"00", -- $00350
          x"06", -- $00351
          x"00", -- $00352
          x"06", -- $00353
          x"06", -- $00354
          x"06", -- $00355
          x"06", -- $00356
          x"3c", -- $00357
          x"00", -- $00358
          x"60", -- $00359
          x"60", -- $0035a
          x"6c", -- $0035b
          x"78", -- $0035c
          x"6c", -- $0035d
          x"66", -- $0035e
          x"00", -- $0035f
          x"00", -- $00360
          x"38", -- $00361
          x"18", -- $00362
          x"18", -- $00363
          x"18", -- $00364
          x"18", -- $00365
          x"3c", -- $00366
          x"00", -- $00367
          x"00", -- $00368
          x"00", -- $00369
          x"66", -- $0036a
          x"7f", -- $0036b
          x"6b", -- $0036c
          x"63", -- $0036d
          x"63", -- $0036e
          x"00", -- $0036f
          x"00", -- $00370
          x"00", -- $00371
          x"7c", -- $00372
          x"66", -- $00373
          x"66", -- $00374
          x"66", -- $00375
          x"66", -- $00376
          x"00", -- $00377
          x"00", -- $00378
          x"00", -- $00379
          x"3c", -- $0037a
          x"66", -- $0037b
          x"66", -- $0037c
          x"66", -- $0037d
          x"3c", -- $0037e
          x"00", -- $0037f
          x"00", -- $00380
          x"00", -- $00381
          x"7c", -- $00382
          x"66", -- $00383
          x"66", -- $00384
          x"7c", -- $00385
          x"60", -- $00386
          x"60", -- $00387
          x"00", -- $00388
          x"00", -- $00389
          x"3e", -- $0038a
          x"66", -- $0038b
          x"66", -- $0038c
          x"3e", -- $0038d
          x"06", -- $0038e
          x"06", -- $0038f
          x"00", -- $00390
          x"00", -- $00391
          x"7c", -- $00392
          x"66", -- $00393
          x"60", -- $00394
          x"60", -- $00395
          x"60", -- $00396
          x"00", -- $00397
          x"00", -- $00398
          x"00", -- $00399
          x"3e", -- $0039a
          x"60", -- $0039b
          x"3c", -- $0039c
          x"06", -- $0039d
          x"7c", -- $0039e
          x"00", -- $0039f
          x"00", -- $003a0
          x"18", -- $003a1
          x"7e", -- $003a2
          x"18", -- $003a3
          x"18", -- $003a4
          x"18", -- $003a5
          x"0e", -- $003a6
          x"00", -- $003a7
          x"00", -- $003a8
          x"00", -- $003a9
          x"66", -- $003aa
          x"66", -- $003ab
          x"66", -- $003ac
          x"66", -- $003ad
          x"3e", -- $003ae
          x"00", -- $003af
          x"00", -- $003b0
          x"00", -- $003b1
          x"66", -- $003b2
          x"66", -- $003b3
          x"66", -- $003b4
          x"3c", -- $003b5
          x"18", -- $003b6
          x"00", -- $003b7
          x"00", -- $003b8
          x"00", -- $003b9
          x"63", -- $003ba
          x"6b", -- $003bb
          x"7f", -- $003bc
          x"3e", -- $003bd
          x"36", -- $003be
          x"00", -- $003bf
          x"00", -- $003c0
          x"00", -- $003c1
          x"66", -- $003c2
          x"3c", -- $003c3
          x"18", -- $003c4
          x"3c", -- $003c5
          x"66", -- $003c6
          x"00", -- $003c7
          x"00", -- $003c8
          x"00", -- $003c9
          x"66", -- $003ca
          x"66", -- $003cb
          x"66", -- $003cc
          x"3e", -- $003cd
          x"0c", -- $003ce
          x"78", -- $003cf
          x"00", -- $003d0
          x"00", -- $003d1
          x"7e", -- $003d2
          x"0c", -- $003d3
          x"18", -- $003d4
          x"30", -- $003d5
          x"7e", -- $003d6
          x"00", -- $003d7
          x"0c", -- $003d8
          x"10", -- $003d9
          x"10", -- $003da
          x"60", -- $003db
          x"10", -- $003dc
          x"10", -- $003dd
          x"0c", -- $003de
          x"00", -- $003df
          x"18", -- $003e0
          x"18", -- $003e1
          x"18", -- $003e2
          x"00", -- $003e3
          x"18", -- $003e4
          x"18", -- $003e5
          x"18", -- $003e6
          x"00", -- $003e7
          x"60", -- $003e8
          x"10", -- $003e9
          x"10", -- $003ea
          x"0c", -- $003eb
          x"10", -- $003ec
          x"10", -- $003ed
          x"60", -- $003ee
          x"00", -- $003ef
          x"00", -- $003f0
          x"32", -- $003f1
          x"4c", -- $003f2
          x"00", -- $003f3
          x"00", -- $003f4
          x"00", -- $003f5
          x"00", -- $003f6
          x"00", -- $003f7
          x"10", -- $003f8
          x"28", -- $003f9
          x"44", -- $003fa
          x"82", -- $003fb
          x"82", -- $003fc
          x"82", -- $003fd
          x"fe", -- $003fe
          x"00", -- $003ff
          x"78", -- $00400
          x"cc", -- $00401
          x"dc", -- $00402
          x"dc", -- $00403
          x"c0", -- $00404
          x"cc", -- $00405
          x"7c", -- $00406
          x"00", -- $00407
          x"78", -- $00408
          x"cc", -- $00409
          x"cc", -- $0040a
          x"fc", -- $0040b
          x"cc", -- $0040c
          x"cc", -- $0040d
          x"cc", -- $0040e
          x"00", -- $0040f
          x"f8", -- $00410
          x"cc", -- $00411
          x"cc", -- $00412
          x"f8", -- $00413
          x"cc", -- $00414
          x"cc", -- $00415
          x"fc", -- $00416
          x"00", -- $00417
          x"78", -- $00418
          x"cc", -- $00419
          x"cc", -- $0041a
          x"c0", -- $0041b
          x"c0", -- $0041c
          x"cc", -- $0041d
          x"7c", -- $0041e
          x"00", -- $0041f
          x"f8", -- $00420
          x"cc", -- $00421
          x"cc", -- $00422
          x"cc", -- $00423
          x"cc", -- $00424
          x"cc", -- $00425
          x"f8", -- $00426
          x"00", -- $00427
          x"fc", -- $00428
          x"cc", -- $00429
          x"c0", -- $0042a
          x"f0", -- $0042b
          x"c0", -- $0042c
          x"cc", -- $0042d
          x"fc", -- $0042e
          x"00", -- $0042f
          x"fc", -- $00430
          x"cc", -- $00431
          x"c0", -- $00432
          x"f0", -- $00433
          x"c0", -- $00434
          x"c0", -- $00435
          x"c0", -- $00436
          x"00", -- $00437
          x"7c", -- $00438
          x"cc", -- $00439
          x"c0", -- $0043a
          x"dc", -- $0043b
          x"cc", -- $0043c
          x"cc", -- $0043d
          x"7c", -- $0043e
          x"00", -- $0043f
          x"cc", -- $00440
          x"cc", -- $00441
          x"cc", -- $00442
          x"fc", -- $00443
          x"cc", -- $00444
          x"cc", -- $00445
          x"cc", -- $00446
          x"00", -- $00447
          x"fc", -- $00448
          x"30", -- $00449
          x"30", -- $0044a
          x"30", -- $0044b
          x"30", -- $0044c
          x"30", -- $0044d
          x"fc", -- $0044e
          x"00", -- $0044f
          x"fc", -- $00450
          x"cc", -- $00451
          x"0c", -- $00452
          x"0c", -- $00453
          x"cc", -- $00454
          x"cc", -- $00455
          x"f8", -- $00456
          x"00", -- $00457
          x"cc", -- $00458
          x"cc", -- $00459
          x"d8", -- $0045a
          x"f0", -- $0045b
          x"d8", -- $0045c
          x"cc", -- $0045d
          x"cc", -- $0045e
          x"00", -- $0045f
          x"c0", -- $00460
          x"c0", -- $00461
          x"c0", -- $00462
          x"c0", -- $00463
          x"c0", -- $00464
          x"cc", -- $00465
          x"fc", -- $00466
          x"00", -- $00467
          x"c6", -- $00468
          x"ee", -- $00469
          x"fe", -- $0046a
          x"fe", -- $0046b
          x"d6", -- $0046c
          x"c6", -- $0046d
          x"c6", -- $0046e
          x"00", -- $0046f
          x"cc", -- $00470
          x"cc", -- $00471
          x"ec", -- $00472
          x"fc", -- $00473
          x"dc", -- $00474
          x"cc", -- $00475
          x"cc", -- $00476
          x"00", -- $00477
          x"78", -- $00478
          x"cc", -- $00479
          x"cc", -- $0047a
          x"cc", -- $0047b
          x"cc", -- $0047c
          x"cc", -- $0047d
          x"7c", -- $0047e
          x"00", -- $0047f
          x"f8", -- $00480
          x"cc", -- $00481
          x"cc", -- $00482
          x"fc", -- $00483
          x"c0", -- $00484
          x"c0", -- $00485
          x"c0", -- $00486
          x"00", -- $00487
          x"78", -- $00488
          x"cc", -- $00489
          x"cc", -- $0048a
          x"cc", -- $0048b
          x"d4", -- $0048c
          x"d8", -- $0048d
          x"6c", -- $0048e
          x"00", -- $0048f
          x"f8", -- $00490
          x"cc", -- $00491
          x"cc", -- $00492
          x"f8", -- $00493
          x"cc", -- $00494
          x"cc", -- $00495
          x"cc", -- $00496
          x"00", -- $00497
          x"7c", -- $00498
          x"c0", -- $00499
          x"e0", -- $0049a
          x"78", -- $0049b
          x"1c", -- $0049c
          x"1c", -- $0049d
          x"f8", -- $0049e
          x"00", -- $0049f
          x"fc", -- $004a0
          x"30", -- $004a1
          x"30", -- $004a2
          x"30", -- $004a3
          x"30", -- $004a4
          x"30", -- $004a5
          x"30", -- $004a6
          x"00", -- $004a7
          x"cc", -- $004a8
          x"cc", -- $004a9
          x"cc", -- $004aa
          x"cc", -- $004ab
          x"cc", -- $004ac
          x"dc", -- $004ad
          x"78", -- $004ae
          x"00", -- $004af
          x"cc", -- $004b0
          x"cc", -- $004b1
          x"cc", -- $004b2
          x"58", -- $004b3
          x"78", -- $004b4
          x"30", -- $004b5
          x"30", -- $004b6
          x"00", -- $004b7
          x"c6", -- $004b8
          x"c6", -- $004b9
          x"d6", -- $004ba
          x"fe", -- $004bb
          x"fe", -- $004bc
          x"ee", -- $004bd
          x"c6", -- $004be
          x"00", -- $004bf
          x"cc", -- $004c0
          x"cc", -- $004c1
          x"78", -- $004c2
          x"30", -- $004c3
          x"78", -- $004c4
          x"cc", -- $004c5
          x"cc", -- $004c6
          x"00", -- $004c7
          x"cc", -- $004c8
          x"cc", -- $004c9
          x"dc", -- $004ca
          x"78", -- $004cb
          x"30", -- $004cc
          x"30", -- $004cd
          x"30", -- $004ce
          x"00", -- $004cf
          x"fc", -- $004d0
          x"cc", -- $004d1
          x"18", -- $004d2
          x"30", -- $004d3
          x"60", -- $004d4
          x"ec", -- $004d5
          x"fc", -- $004d6
          x"00", -- $004d7
          x"78", -- $004d8
          x"60", -- $004d9
          x"60", -- $004da
          x"60", -- $004db
          x"60", -- $004dc
          x"60", -- $004dd
          x"78", -- $004de
          x"00", -- $004df
          x"78", -- $004e0
          x"cc", -- $004e1
          x"c0", -- $004e2
          x"f0", -- $004e3
          x"60", -- $004e4
          x"60", -- $004e5
          x"fc", -- $004e6
          x"00", -- $004e7
          x"78", -- $004e8
          x"18", -- $004e9
          x"18", -- $004ea
          x"18", -- $004eb
          x"18", -- $004ec
          x"18", -- $004ed
          x"78", -- $004ee
          x"00", -- $004ef
          x"10", -- $004f0
          x"38", -- $004f1
          x"7c", -- $004f2
          x"38", -- $004f3
          x"38", -- $004f4
          x"38", -- $004f5
          x"38", -- $004f6
          x"00", -- $004f7
          x"00", -- $004f8
          x"20", -- $004f9
          x"7e", -- $004fa
          x"fe", -- $004fb
          x"7e", -- $004fc
          x"20", -- $004fd
          x"00", -- $004fe
          x"00", -- $004ff
          x"00", -- $00500
          x"00", -- $00501
          x"00", -- $00502
          x"00", -- $00503
          x"00", -- $00504
          x"00", -- $00505
          x"00", -- $00506
          x"00", -- $00507
          x"00", -- $00508
          x"00", -- $00509
          x"00", -- $0050a
          x"00", -- $0050b
          x"00", -- $0050c
          x"00", -- $0050d
          x"00", -- $0050e
          x"00", -- $0050f
          x"00", -- $00510
          x"00", -- $00511
          x"00", -- $00512
          x"00", -- $00513
          x"00", -- $00514
          x"00", -- $00515
          x"00", -- $00516
          x"00", -- $00517
          x"00", -- $00518
          x"00", -- $00519
          x"00", -- $0051a
          x"00", -- $0051b
          x"00", -- $0051c
          x"00", -- $0051d
          x"00", -- $0051e
          x"00", -- $0051f
          x"00", -- $00520
          x"00", -- $00521
          x"00", -- $00522
          x"00", -- $00523
          x"00", -- $00524
          x"00", -- $00525
          x"00", -- $00526
          x"00", -- $00527
          x"00", -- $00528
          x"00", -- $00529
          x"00", -- $0052a
          x"00", -- $0052b
          x"00", -- $0052c
          x"00", -- $0052d
          x"00", -- $0052e
          x"00", -- $0052f
          x"00", -- $00530
          x"00", -- $00531
          x"00", -- $00532
          x"00", -- $00533
          x"00", -- $00534
          x"00", -- $00535
          x"00", -- $00536
          x"00", -- $00537
          x"00", -- $00538
          x"00", -- $00539
          x"00", -- $0053a
          x"00", -- $0053b
          x"00", -- $0053c
          x"00", -- $0053d
          x"00", -- $0053e
          x"00", -- $0053f
          x"00", -- $00540
          x"00", -- $00541
          x"00", -- $00542
          x"00", -- $00543
          x"00", -- $00544
          x"00", -- $00545
          x"00", -- $00546
          x"00", -- $00547
          x"00", -- $00548
          x"00", -- $00549
          x"00", -- $0054a
          x"00", -- $0054b
          x"00", -- $0054c
          x"00", -- $0054d
          x"00", -- $0054e
          x"00", -- $0054f
          x"00", -- $00550
          x"00", -- $00551
          x"00", -- $00552
          x"00", -- $00553
          x"00", -- $00554
          x"00", -- $00555
          x"00", -- $00556
          x"00", -- $00557
          x"00", -- $00558
          x"00", -- $00559
          x"00", -- $0055a
          x"00", -- $0055b
          x"00", -- $0055c
          x"00", -- $0055d
          x"00", -- $0055e
          x"00", -- $0055f
          x"00", -- $00560
          x"00", -- $00561
          x"00", -- $00562
          x"00", -- $00563
          x"00", -- $00564
          x"00", -- $00565
          x"00", -- $00566
          x"00", -- $00567
          x"00", -- $00568
          x"00", -- $00569
          x"00", -- $0056a
          x"00", -- $0056b
          x"00", -- $0056c
          x"00", -- $0056d
          x"00", -- $0056e
          x"00", -- $0056f
          x"00", -- $00570
          x"00", -- $00571
          x"00", -- $00572
          x"00", -- $00573
          x"00", -- $00574
          x"00", -- $00575
          x"00", -- $00576
          x"00", -- $00577
          x"00", -- $00578
          x"00", -- $00579
          x"00", -- $0057a
          x"00", -- $0057b
          x"00", -- $0057c
          x"00", -- $0057d
          x"00", -- $0057e
          x"00", -- $0057f
          x"00", -- $00580
          x"00", -- $00581
          x"00", -- $00582
          x"00", -- $00583
          x"00", -- $00584
          x"00", -- $00585
          x"00", -- $00586
          x"00", -- $00587
          x"00", -- $00588
          x"00", -- $00589
          x"00", -- $0058a
          x"00", -- $0058b
          x"00", -- $0058c
          x"00", -- $0058d
          x"00", -- $0058e
          x"00", -- $0058f
          x"00", -- $00590
          x"00", -- $00591
          x"00", -- $00592
          x"00", -- $00593
          x"00", -- $00594
          x"00", -- $00595
          x"00", -- $00596
          x"00", -- $00597
          x"00", -- $00598
          x"00", -- $00599
          x"00", -- $0059a
          x"00", -- $0059b
          x"00", -- $0059c
          x"00", -- $0059d
          x"00", -- $0059e
          x"00", -- $0059f
          x"00", -- $005a0
          x"00", -- $005a1
          x"00", -- $005a2
          x"00", -- $005a3
          x"00", -- $005a4
          x"00", -- $005a5
          x"00", -- $005a6
          x"00", -- $005a7
          x"00", -- $005a8
          x"00", -- $005a9
          x"00", -- $005aa
          x"00", -- $005ab
          x"00", -- $005ac
          x"00", -- $005ad
          x"00", -- $005ae
          x"00", -- $005af
          x"00", -- $005b0
          x"00", -- $005b1
          x"00", -- $005b2
          x"00", -- $005b3
          x"00", -- $005b4
          x"00", -- $005b5
          x"00", -- $005b6
          x"00", -- $005b7
          x"00", -- $005b8
          x"00", -- $005b9
          x"00", -- $005ba
          x"00", -- $005bb
          x"00", -- $005bc
          x"00", -- $005bd
          x"00", -- $005be
          x"00", -- $005bf
          x"00", -- $005c0
          x"00", -- $005c1
          x"00", -- $005c2
          x"00", -- $005c3
          x"00", -- $005c4
          x"00", -- $005c5
          x"00", -- $005c6
          x"00", -- $005c7
          x"00", -- $005c8
          x"00", -- $005c9
          x"00", -- $005ca
          x"00", -- $005cb
          x"00", -- $005cc
          x"00", -- $005cd
          x"00", -- $005ce
          x"00", -- $005cf
          x"00", -- $005d0
          x"00", -- $005d1
          x"00", -- $005d2
          x"00", -- $005d3
          x"00", -- $005d4
          x"00", -- $005d5
          x"00", -- $005d6
          x"00", -- $005d7
          x"00", -- $005d8
          x"00", -- $005d9
          x"00", -- $005da
          x"00", -- $005db
          x"00", -- $005dc
          x"00", -- $005dd
          x"00", -- $005de
          x"00", -- $005df
          x"00", -- $005e0
          x"00", -- $005e1
          x"00", -- $005e2
          x"00", -- $005e3
          x"00", -- $005e4
          x"00", -- $005e5
          x"00", -- $005e6
          x"00", -- $005e7
          x"00", -- $005e8
          x"00", -- $005e9
          x"00", -- $005ea
          x"00", -- $005eb
          x"00", -- $005ec
          x"00", -- $005ed
          x"00", -- $005ee
          x"00", -- $005ef
          x"00", -- $005f0
          x"00", -- $005f1
          x"00", -- $005f2
          x"00", -- $005f3
          x"00", -- $005f4
          x"00", -- $005f5
          x"00", -- $005f6
          x"00", -- $005f7
          x"00", -- $005f8
          x"00", -- $005f9
          x"00", -- $005fa
          x"00", -- $005fb
          x"00", -- $005fc
          x"00", -- $005fd
          x"00", -- $005fe
          x"00", -- $005ff
          x"00", -- $00600
          x"00", -- $00601
          x"00", -- $00602
          x"00", -- $00603
          x"00", -- $00604
          x"00", -- $00605
          x"00", -- $00606
          x"00", -- $00607
          x"00", -- $00608
          x"00", -- $00609
          x"00", -- $0060a
          x"00", -- $0060b
          x"00", -- $0060c
          x"00", -- $0060d
          x"00", -- $0060e
          x"00", -- $0060f
          x"00", -- $00610
          x"00", -- $00611
          x"00", -- $00612
          x"00", -- $00613
          x"00", -- $00614
          x"00", -- $00615
          x"00", -- $00616
          x"00", -- $00617
          x"00", -- $00618
          x"00", -- $00619
          x"00", -- $0061a
          x"00", -- $0061b
          x"00", -- $0061c
          x"00", -- $0061d
          x"00", -- $0061e
          x"00", -- $0061f
          x"00", -- $00620
          x"00", -- $00621
          x"00", -- $00622
          x"00", -- $00623
          x"00", -- $00624
          x"00", -- $00625
          x"00", -- $00626
          x"00", -- $00627
          x"00", -- $00628
          x"00", -- $00629
          x"00", -- $0062a
          x"00", -- $0062b
          x"00", -- $0062c
          x"00", -- $0062d
          x"00", -- $0062e
          x"00", -- $0062f
          x"00", -- $00630
          x"00", -- $00631
          x"00", -- $00632
          x"00", -- $00633
          x"00", -- $00634
          x"00", -- $00635
          x"00", -- $00636
          x"00", -- $00637
          x"00", -- $00638
          x"00", -- $00639
          x"00", -- $0063a
          x"00", -- $0063b
          x"00", -- $0063c
          x"00", -- $0063d
          x"00", -- $0063e
          x"00", -- $0063f
          x"00", -- $00640
          x"00", -- $00641
          x"00", -- $00642
          x"00", -- $00643
          x"00", -- $00644
          x"00", -- $00645
          x"00", -- $00646
          x"00", -- $00647
          x"00", -- $00648
          x"00", -- $00649
          x"00", -- $0064a
          x"00", -- $0064b
          x"00", -- $0064c
          x"00", -- $0064d
          x"00", -- $0064e
          x"00", -- $0064f
          x"00", -- $00650
          x"00", -- $00651
          x"00", -- $00652
          x"00", -- $00653
          x"00", -- $00654
          x"00", -- $00655
          x"00", -- $00656
          x"00", -- $00657
          x"00", -- $00658
          x"00", -- $00659
          x"00", -- $0065a
          x"00", -- $0065b
          x"00", -- $0065c
          x"00", -- $0065d
          x"00", -- $0065e
          x"00", -- $0065f
          x"00", -- $00660
          x"00", -- $00661
          x"00", -- $00662
          x"00", -- $00663
          x"00", -- $00664
          x"00", -- $00665
          x"00", -- $00666
          x"00", -- $00667
          x"00", -- $00668
          x"00", -- $00669
          x"00", -- $0066a
          x"00", -- $0066b
          x"00", -- $0066c
          x"00", -- $0066d
          x"00", -- $0066e
          x"00", -- $0066f
          x"00", -- $00670
          x"00", -- $00671
          x"00", -- $00672
          x"00", -- $00673
          x"00", -- $00674
          x"00", -- $00675
          x"00", -- $00676
          x"00", -- $00677
          x"00", -- $00678
          x"00", -- $00679
          x"00", -- $0067a
          x"00", -- $0067b
          x"00", -- $0067c
          x"00", -- $0067d
          x"00", -- $0067e
          x"00", -- $0067f
          x"00", -- $00680
          x"00", -- $00681
          x"00", -- $00682
          x"00", -- $00683
          x"00", -- $00684
          x"00", -- $00685
          x"00", -- $00686
          x"00", -- $00687
          x"00", -- $00688
          x"00", -- $00689
          x"00", -- $0068a
          x"00", -- $0068b
          x"00", -- $0068c
          x"00", -- $0068d
          x"00", -- $0068e
          x"00", -- $0068f
          x"00", -- $00690
          x"00", -- $00691
          x"00", -- $00692
          x"00", -- $00693
          x"00", -- $00694
          x"00", -- $00695
          x"00", -- $00696
          x"00", -- $00697
          x"00", -- $00698
          x"00", -- $00699
          x"00", -- $0069a
          x"00", -- $0069b
          x"00", -- $0069c
          x"00", -- $0069d
          x"00", -- $0069e
          x"00", -- $0069f
          x"00", -- $006a0
          x"00", -- $006a1
          x"00", -- $006a2
          x"00", -- $006a3
          x"00", -- $006a4
          x"00", -- $006a5
          x"00", -- $006a6
          x"00", -- $006a7
          x"00", -- $006a8
          x"00", -- $006a9
          x"00", -- $006aa
          x"00", -- $006ab
          x"00", -- $006ac
          x"00", -- $006ad
          x"00", -- $006ae
          x"00", -- $006af
          x"00", -- $006b0
          x"00", -- $006b1
          x"00", -- $006b2
          x"00", -- $006b3
          x"00", -- $006b4
          x"00", -- $006b5
          x"00", -- $006b6
          x"00", -- $006b7
          x"00", -- $006b8
          x"00", -- $006b9
          x"00", -- $006ba
          x"00", -- $006bb
          x"00", -- $006bc
          x"00", -- $006bd
          x"00", -- $006be
          x"00", -- $006bf
          x"00", -- $006c0
          x"00", -- $006c1
          x"00", -- $006c2
          x"00", -- $006c3
          x"00", -- $006c4
          x"00", -- $006c5
          x"00", -- $006c6
          x"00", -- $006c7
          x"00", -- $006c8
          x"00", -- $006c9
          x"00", -- $006ca
          x"00", -- $006cb
          x"00", -- $006cc
          x"00", -- $006cd
          x"00", -- $006ce
          x"00", -- $006cf
          x"00", -- $006d0
          x"00", -- $006d1
          x"00", -- $006d2
          x"00", -- $006d3
          x"00", -- $006d4
          x"00", -- $006d5
          x"00", -- $006d6
          x"00", -- $006d7
          x"00", -- $006d8
          x"00", -- $006d9
          x"00", -- $006da
          x"00", -- $006db
          x"00", -- $006dc
          x"00", -- $006dd
          x"00", -- $006de
          x"00", -- $006df
          x"00", -- $006e0
          x"00", -- $006e1
          x"00", -- $006e2
          x"00", -- $006e3
          x"00", -- $006e4
          x"00", -- $006e5
          x"00", -- $006e6
          x"00", -- $006e7
          x"00", -- $006e8
          x"00", -- $006e9
          x"00", -- $006ea
          x"00", -- $006eb
          x"00", -- $006ec
          x"00", -- $006ed
          x"00", -- $006ee
          x"00", -- $006ef
          x"00", -- $006f0
          x"00", -- $006f1
          x"00", -- $006f2
          x"00", -- $006f3
          x"00", -- $006f4
          x"00", -- $006f5
          x"00", -- $006f6
          x"00", -- $006f7
          x"00", -- $006f8
          x"00", -- $006f9
          x"00", -- $006fa
          x"00", -- $006fb
          x"00", -- $006fc
          x"00", -- $006fd
          x"00", -- $006fe
          x"00", -- $006ff
          x"00", -- $00700
          x"00", -- $00701
          x"00", -- $00702
          x"00", -- $00703
          x"00", -- $00704
          x"00", -- $00705
          x"00", -- $00706
          x"00", -- $00707
          x"00", -- $00708
          x"00", -- $00709
          x"00", -- $0070a
          x"00", -- $0070b
          x"00", -- $0070c
          x"00", -- $0070d
          x"00", -- $0070e
          x"00", -- $0070f
          x"00", -- $00710
          x"00", -- $00711
          x"00", -- $00712
          x"00", -- $00713
          x"00", -- $00714
          x"00", -- $00715
          x"00", -- $00716
          x"00", -- $00717
          x"00", -- $00718
          x"00", -- $00719
          x"00", -- $0071a
          x"00", -- $0071b
          x"00", -- $0071c
          x"00", -- $0071d
          x"00", -- $0071e
          x"00", -- $0071f
          x"00", -- $00720
          x"00", -- $00721
          x"00", -- $00722
          x"00", -- $00723
          x"00", -- $00724
          x"00", -- $00725
          x"00", -- $00726
          x"00", -- $00727
          x"00", -- $00728
          x"00", -- $00729
          x"00", -- $0072a
          x"00", -- $0072b
          x"00", -- $0072c
          x"00", -- $0072d
          x"00", -- $0072e
          x"00", -- $0072f
          x"00", -- $00730
          x"00", -- $00731
          x"00", -- $00732
          x"00", -- $00733
          x"00", -- $00734
          x"00", -- $00735
          x"00", -- $00736
          x"00", -- $00737
          x"00", -- $00738
          x"00", -- $00739
          x"00", -- $0073a
          x"00", -- $0073b
          x"00", -- $0073c
          x"00", -- $0073d
          x"00", -- $0073e
          x"00", -- $0073f
          x"00", -- $00740
          x"00", -- $00741
          x"00", -- $00742
          x"00", -- $00743
          x"00", -- $00744
          x"00", -- $00745
          x"00", -- $00746
          x"00", -- $00747
          x"00", -- $00748
          x"00", -- $00749
          x"00", -- $0074a
          x"00", -- $0074b
          x"00", -- $0074c
          x"00", -- $0074d
          x"00", -- $0074e
          x"00", -- $0074f
          x"00", -- $00750
          x"00", -- $00751
          x"00", -- $00752
          x"00", -- $00753
          x"00", -- $00754
          x"00", -- $00755
          x"00", -- $00756
          x"00", -- $00757
          x"00", -- $00758
          x"00", -- $00759
          x"00", -- $0075a
          x"00", -- $0075b
          x"00", -- $0075c
          x"00", -- $0075d
          x"00", -- $0075e
          x"00", -- $0075f
          x"00", -- $00760
          x"00", -- $00761
          x"00", -- $00762
          x"00", -- $00763
          x"00", -- $00764
          x"00", -- $00765
          x"00", -- $00766
          x"00", -- $00767
          x"00", -- $00768
          x"00", -- $00769
          x"00", -- $0076a
          x"00", -- $0076b
          x"00", -- $0076c
          x"00", -- $0076d
          x"00", -- $0076e
          x"00", -- $0076f
          x"00", -- $00770
          x"00", -- $00771
          x"00", -- $00772
          x"00", -- $00773
          x"00", -- $00774
          x"00", -- $00775
          x"00", -- $00776
          x"00", -- $00777
          x"00", -- $00778
          x"00", -- $00779
          x"00", -- $0077a
          x"00", -- $0077b
          x"00", -- $0077c
          x"00", -- $0077d
          x"00", -- $0077e
          x"00", -- $0077f
          x"00", -- $00780
          x"00", -- $00781
          x"00", -- $00782
          x"00", -- $00783
          x"00", -- $00784
          x"00", -- $00785
          x"00", -- $00786
          x"00", -- $00787
          x"00", -- $00788
          x"00", -- $00789
          x"00", -- $0078a
          x"00", -- $0078b
          x"00", -- $0078c
          x"00", -- $0078d
          x"00", -- $0078e
          x"00", -- $0078f
          x"00", -- $00790
          x"00", -- $00791
          x"00", -- $00792
          x"00", -- $00793
          x"00", -- $00794
          x"00", -- $00795
          x"00", -- $00796
          x"00", -- $00797
          x"00", -- $00798
          x"00", -- $00799
          x"00", -- $0079a
          x"00", -- $0079b
          x"00", -- $0079c
          x"00", -- $0079d
          x"00", -- $0079e
          x"00", -- $0079f
          x"00", -- $007a0
          x"00", -- $007a1
          x"00", -- $007a2
          x"00", -- $007a3
          x"00", -- $007a4
          x"00", -- $007a5
          x"00", -- $007a6
          x"00", -- $007a7
          x"00", -- $007a8
          x"00", -- $007a9
          x"00", -- $007aa
          x"00", -- $007ab
          x"00", -- $007ac
          x"00", -- $007ad
          x"00", -- $007ae
          x"00", -- $007af
          x"00", -- $007b0
          x"00", -- $007b1
          x"00", -- $007b2
          x"00", -- $007b3
          x"00", -- $007b4
          x"00", -- $007b5
          x"00", -- $007b6
          x"00", -- $007b7
          x"00", -- $007b8
          x"00", -- $007b9
          x"00", -- $007ba
          x"00", -- $007bb
          x"00", -- $007bc
          x"00", -- $007bd
          x"00", -- $007be
          x"00", -- $007bf
          x"0f", -- $007c0
          x"0f", -- $007c1
          x"0f", -- $007c2
          x"ff", -- $007c3
          x"fe", -- $007c4
          x"fc", -- $007c5
          x"00", -- $007c6
          x"00", -- $007c7
          x"80", -- $007c8
          x"c0", -- $007c9
          x"e0", -- $007ca
          x"80", -- $007cb
          x"80", -- $007cc
          x"80", -- $007cd
          x"80", -- $007ce
          x"80", -- $007cf
          x"f0", -- $007d0
          x"f0", -- $007d1
          x"f0", -- $007d2
          x"ff", -- $007d3
          x"7f", -- $007d4
          x"3f", -- $007d5
          x"00", -- $007d6
          x"00", -- $007d7
          x"01", -- $007d8
          x"03", -- $007d9
          x"07", -- $007da
          x"01", -- $007db
          x"01", -- $007dc
          x"01", -- $007dd
          x"01", -- $007de
          x"01", -- $007df
          x"01", -- $007e0
          x"01", -- $007e1
          x"01", -- $007e2
          x"01", -- $007e3
          x"01", -- $007e4
          x"07", -- $007e5
          x"03", -- $007e6
          x"01", -- $007e7
          x"00", -- $007e8
          x"00", -- $007e9
          x"3f", -- $007ea
          x"7f", -- $007eb
          x"ff", -- $007ec
          x"f0", -- $007ed
          x"f0", -- $007ee
          x"f0", -- $007ef
          x"80", -- $007f0
          x"80", -- $007f1
          x"80", -- $007f2
          x"80", -- $007f3
          x"80", -- $007f4
          x"e0", -- $007f5
          x"c0", -- $007f6
          x"80", -- $007f7
          x"00", -- $007f8
          x"00", -- $007f9
          x"fc", -- $007fa
          x"fe", -- $007fb
          x"ff", -- $007fc
          x"0f", -- $007fd
          x"0f", -- $007fe
          x"0f", -- $007ff
          x"3f", -- $00800
          x"7f", -- $00801
          x"47", -- $00802
          x"42", -- $00803
          x"50", -- $00804
          x"40", -- $00805
          x"7f", -- $00806
          x"04", -- $00807
          x"05", -- $00808
          x"06", -- $00809
          x"03", -- $0080a
          x"7f", -- $0080b
          x"44", -- $0080c
          x"45", -- $0080d
          x"46", -- $0080e
          x"43", -- $0080f
          x"39", -- $00810
          x"38", -- $00811
          x"3b", -- $00812
          x"08", -- $00813
          x"0b", -- $00814
          x"10", -- $00815
          x"13", -- $00816
          x"18", -- $00817
          x"1b", -- $00818
          x"20", -- $00819
          x"23", -- $0081a
          x"28", -- $0081b
          x"2b", -- $0081c
          x"30", -- $0081d
          x"33", -- $0081e
          x"00", -- $0081f
          x"c1", -- $00820
          x"3e", -- $00821
          x"09", -- $00822
          x"0e", -- $00823
          x"11", -- $00824
          x"16", -- $00825
          x"19", -- $00826
          x"1e", -- $00827
          x"21", -- $00828
          x"26", -- $00829
          x"29", -- $0082a
          x"2e", -- $0082b
          x"31", -- $0082c
          x"36", -- $0082d
          x"d1", -- $0082e
          x"7f", -- $0082f
          x"3a", -- $00830
          x"0f", -- $00831
          x"0a", -- $00832
          x"0d", -- $00833
          x"12", -- $00834
          x"15", -- $00835
          x"1a", -- $00836
          x"1d", -- $00837
          x"22", -- $00838
          x"25", -- $00839
          x"2a", -- $0083a
          x"2d", -- $0083b
          x"32", -- $0083c
          x"35", -- $0083d
          x"01", -- $0083e
          x"01", -- $0083f
          x"3d", -- $00840
          x"8f", -- $00841
          x"0c", -- $00842
          x"17", -- $00843
          x"14", -- $00844
          x"1f", -- $00845
          x"1c", -- $00846
          x"27", -- $00847
          x"24", -- $00848
          x"2f", -- $00849
          x"2c", -- $0084a
          x"37", -- $0084b
          x"b4", -- $0084c
          x"52", -- $0084d
          x"7e", -- $0084e
          x"7e", -- $0084f
          x"7e", -- $00850
          x"7e", -- $00851
          x"7e", -- $00852
          x"3c", -- $00853
          x"3c", -- $00854
          x"3c", -- $00855
          x"3c", -- $00856
          x"3c", -- $00857
          x"3c", -- $00858
          x"3c", -- $00859
          x"3c", -- $0085a
          x"3c", -- $0085b
          x"7e", -- $0085c
          x"53", -- $0085d
          x"07", -- $0085e
          x"02", -- $0085f
          x"7f", -- $00860
          x"7f", -- $00861
          x"7f", -- $00862
          x"7e", -- $00863
          x"7e", -- $00864
          x"7e", -- $00865
          x"7e", -- $00866
          x"7e", -- $00867
          x"7e", -- $00868
          x"7e", -- $00869
          x"7e", -- $0086a
          x"7e", -- $0086b
          x"7f", -- $0086c
          x"7e", -- $0086d
          x"7e", -- $0086e
          x"7e", -- $0086f
          x"7f", -- $00870
          x"7f", -- $00871
          x"7f", -- $00872
          x"7f", -- $00873
          x"7f", -- $00874
          x"7f", -- $00875
          x"7f", -- $00876
          x"7f", -- $00877
          x"7f", -- $00878
          x"7f", -- $00879
          x"7f", -- $0087a
          x"7f", -- $0087b
          x"7f", -- $0087c
          x"7f", -- $0087d
          x"7f", -- $0087e
          x"7f", -- $0087f
          x"7f", -- $00880
          x"38", -- $00881
          x"3b", -- $00882
          x"08", -- $00883
          x"7f", -- $00884
          x"21", -- $00885
          x"7f", -- $00886
          x"04", -- $00887
          x"7f", -- $00888
          x"7f", -- $00889
          x"7f", -- $0088a
          x"7f", -- $0088b
          x"7f", -- $0088c
          x"7f", -- $0088d
          x"7f", -- $0088e
          x"7f", -- $0088f
          x"7f", -- $00890
          x"0b", -- $00891
          x"10", -- $00892
          x"13", -- $00893
          x"7f", -- $00894
          x"7e", -- $00895
          x"7f", -- $00896
          x"05", -- $00897
          x"7f", -- $00898
          x"7f", -- $00899
          x"7f", -- $0089a
          x"7f", -- $0089b
          x"7f", -- $0089c
          x"7f", -- $0089d
          x"7f", -- $0089e
          x"7f", -- $0089f
          x"7f", -- $008a0
          x"18", -- $008a1
          x"1b", -- $008a2
          x"20", -- $008a3
          x"7f", -- $008a4
          x"7f", -- $008a5
          x"7f", -- $008a6
          x"06", -- $008a7
          x"7f", -- $008a8
          x"7f", -- $008a9
          x"7f", -- $008aa
          x"7f", -- $008ab
          x"7f", -- $008ac
          x"7f", -- $008ad
          x"7f", -- $008ae
          x"7f", -- $008af
          x"7f", -- $008b0
          x"37", -- $008b1
          x"23", -- $008b2
          x"31", -- $008b3
          x"7f", -- $008b4
          x"27", -- $008b5
          x"7f", -- $008b6
          x"03", -- $008b7
          x"7f", -- $008b8
          x"7f", -- $008b9
          x"7f", -- $008ba
          x"7f", -- $008bb
          x"7f", -- $008bc
          x"7f", -- $008bd
          x"7f", -- $008be
          x"7f", -- $008bf
          x"7f", -- $008c0
          x"7e", -- $008c1
          x"7e", -- $008c2
          x"7e", -- $008c3
          x"7f", -- $008c4
          x"7e", -- $008c5
          x"7f", -- $008c6
          x"7e", -- $008c7
          x"7f", -- $008c8
          x"7f", -- $008c9
          x"7f", -- $008ca
          x"7f", -- $008cb
          x"7f", -- $008cc
          x"7f", -- $008cd
          x"7f", -- $008ce
          x"7f", -- $008cf
          x"7f", -- $008d0
          x"7f", -- $008d1
          x"7f", -- $008d2
          x"7f", -- $008d3
          x"7f", -- $008d4
          x"7f", -- $008d5
          x"7f", -- $008d6
          x"7f", -- $008d7
          x"7f", -- $008d8
          x"7f", -- $008d9
          x"7f", -- $008da
          x"7f", -- $008db
          x"7f", -- $008dc
          x"7f", -- $008dd
          x"7f", -- $008de
          x"7f", -- $008df
          x"00", -- $008e0
          x"00", -- $008e1
          x"00", -- $008e2
          x"00", -- $008e3
          x"00", -- $008e4
          x"00", -- $008e5
          x"00", -- $008e6
          x"00", -- $008e7
          x"00", -- $008e8
          x"00", -- $008e9
          x"00", -- $008ea
          x"00", -- $008eb
          x"00", -- $008ec
          x"00", -- $008ed
          x"00", -- $008ee
          x"00", -- $008ef
          x"00", -- $008f0
          x"00", -- $008f1
          x"00", -- $008f2
          x"00", -- $008f3
          x"00", -- $008f4
          x"00", -- $008f5
          x"00", -- $008f6
          x"00", -- $008f7
          x"00", -- $008f8
          x"00", -- $008f9
          x"00", -- $008fa
          x"00", -- $008fb
          x"00", -- $008fc
          x"00", -- $008fd
          x"00", -- $008fe
          x"00", -- $008ff
          x"0a", -- $00900
          x"52", -- $00901
          x"55", -- $00902
          x"4e", -- $00903
          x"95", -- $00904
          x"45", -- $00905
          x"53", -- $00906
          x"43", -- $00907
          x"90", -- $00908
          x"41", -- $00909
          x"4c", -- $0090a
          x"54", -- $0090b
          x"90", -- $0090c
          x"41", -- $0090d
          x"53", -- $0090e
          x"43", -- $0090f
          x"91", -- $00910
          x"4e", -- $00911
          x"4f", -- $00912
          x"96", -- $00913
          x"46", -- $00914
          x"31", -- $00915
          x"91", -- $00916
          x"46", -- $00917
          x"33", -- $00918
          x"91", -- $00919
          x"46", -- $0091a
          x"35", -- $0091b
          x"91", -- $0091c
          x"46", -- $0091d
          x"37", -- $0091e
          x"95", -- $0091f
          x"46", -- $00920
          x"39", -- $00921
          x"91", -- $00922
          x"46", -- $00923
          x"31", -- $00924
          x"31", -- $00925
          x"90", -- $00926
          x"46", -- $00927
          x"31", -- $00928
          x"33", -- $00929
          x"90", -- $0092a
          x"48", -- $0092b
          x"45", -- $0092c
          x"4c", -- $0092d
          x"50", -- $0092e
          x"0a", -- $0092f
          x"53", -- $00930
          x"54", -- $00931
          x"4f", -- $00932
          x"50", -- $00933
          x"9e", -- $00934
          x"44", -- $00935
          x"49", -- $00936
          x"4e", -- $00937
          x"90", -- $00938
          x"53", -- $00939
          x"43", -- $0093a
          x"52", -- $0093b
          x"4c", -- $0093c
          x"95", -- $0093d
          x"46", -- $0093e
          x"32", -- $0093f
          x"91", -- $00940
          x"46", -- $00941
          x"34", -- $00942
          x"91", -- $00943
          x"46", -- $00944
          x"36", -- $00945
          x"91", -- $00946
          x"46", -- $00947
          x"38", -- $00948
          x"95", -- $00949
          x"46", -- $0094a
          x"31", -- $0094b
          x"30", -- $0094c
          x"90", -- $0094d
          x"46", -- $0094e
          x"31", -- $0094f
          x"32", -- $00950
          x"90", -- $00951
          x"46", -- $00952
          x"31", -- $00953
          x"34", -- $00954
          x"0a", -- $00955
          x"0a", -- $00956
          x"20", -- $00957
          x"7e", -- $00958
          x"92", -- $00959
          x"21", -- $0095a
          x"92", -- $0095b
          x"22", -- $0095c
          x"92", -- $0095d
          x"23", -- $0095e
          x"92", -- $0095f
          x"24", -- $00960
          x"92", -- $00961
          x"25", -- $00962
          x"92", -- $00963
          x"26", -- $00964
          x"92", -- $00965
          x"27", -- $00966
          x"92", -- $00967
          x"28", -- $00968
          x"92", -- $00969
          x"29", -- $0096a
          x"92", -- $0096b
          x"60", -- $0096c
          x"9f", -- $0096d
          x"20", -- $0096e
          x"43", -- $0096f
          x"4c", -- $00970
          x"52", -- $00971
          x"90", -- $00972
          x"49", -- $00973
          x"4e", -- $00974
          x"53", -- $00975
          x"54", -- $00976
          x"0a", -- $00977
          x"20", -- $00978
          x"5f", -- $00979
          x"92", -- $0097a
          x"31", -- $0097b
          x"92", -- $0097c
          x"32", -- $0097d
          x"92", -- $0097e
          x"33", -- $0097f
          x"92", -- $00980
          x"34", -- $00981
          x"92", -- $00982
          x"35", -- $00983
          x"92", -- $00984
          x"36", -- $00985
          x"92", -- $00986
          x"37", -- $00987
          x"92", -- $00988
          x"38", -- $00989
          x"92", -- $0098a
          x"39", -- $0098b
          x"92", -- $0098c
          x"30", -- $0098d
          x"92", -- $0098e
          x"2b", -- $0098f
          x"92", -- $00990
          x"2d", -- $00991
          x"91", -- $00992
          x"47", -- $00993
          x"42", -- $00994
          x"50", -- $00995
          x"90", -- $00996
          x"48", -- $00997
          x"4f", -- $00998
          x"4d", -- $00999
          x"45", -- $0099a
          x"20", -- $0099b
          x"44", -- $0099c
          x"45", -- $0099d
          x"4c", -- $0099e
          x"0a", -- $0099f
          x"0a", -- $009a0
          x"54", -- $009a1
          x"41", -- $009a2
          x"42", -- $009a3
          x"9f", -- $009a4
          x"9f", -- $009a5
          x"9f", -- $009a6
          x"9d", -- $009a7
          x"50", -- $009a8
          x"49", -- $009a9
          x"0a", -- $009aa
          x"97", -- $009ab
          x"51", -- $009ac
          x"92", -- $009ad
          x"57", -- $009ae
          x"92", -- $009af
          x"45", -- $009b0
          x"92", -- $009b1
          x"52", -- $009b2
          x"92", -- $009b3
          x"54", -- $009b4
          x"92", -- $009b5
          x"59", -- $009b6
          x"92", -- $009b7
          x"55", -- $009b8
          x"92", -- $009b9
          x"49", -- $009ba
          x"92", -- $009bb
          x"4f", -- $009bc
          x"92", -- $009bd
          x"50", -- $009be
          x"92", -- $009bf
          x"40", -- $009c0
          x"92", -- $009c1
          x"2a", -- $009c2
          x"92", -- $009c3
          x"7e", -- $009c4
          x"5e", -- $009c5
          x"90", -- $009c6
          x"52", -- $009c7
          x"45", -- $009c8
          x"53", -- $009c9
          x"54", -- $009ca
          x"4f", -- $009cb
          x"52", -- $009cc
          x"45", -- $009cd
          x"0a", -- $009ce
          x"0a", -- $009cf
          x"43", -- $009d0
          x"54", -- $009d1
          x"52", -- $009d2
          x"4c", -- $009d3
          x"20", -- $009d4
          x"53", -- $009d5
          x"48", -- $009d6
          x"46", -- $009d7
          x"54", -- $009d8
          x"9f", -- $009d9
          x"9f", -- $009da
          x"9b", -- $009db
          x"5b", -- $009dc
          x"92", -- $009dd
          x"5d", -- $009de
          x"0a", -- $009df
          x"93", -- $009e0
          x"4c", -- $009e1
          x"4f", -- $009e2
          x"43", -- $009e3
          x"4b", -- $009e4
          x"90", -- $009e5
          x"41", -- $009e6
          x"92", -- $009e7
          x"53", -- $009e8
          x"92", -- $009e9
          x"44", -- $009ea
          x"92", -- $009eb
          x"46", -- $009ec
          x"92", -- $009ed
          x"47", -- $009ee
          x"92", -- $009ef
          x"48", -- $009f0
          x"92", -- $009f1
          x"4a", -- $009f2
          x"92", -- $009f3
          x"4b", -- $009f4
          x"92", -- $009f5
          x"4c", -- $009f6
          x"92", -- $009f7
          x"7b", -- $009f8
          x"3a", -- $009f9
          x"91", -- $009fa
          x"7d", -- $009fb
          x"3b", -- $009fc
          x"91", -- $009fd
          x"3d", -- $009fe
          x"93", -- $009ff
          x"52", -- $00a00
          x"45", -- $00a01
          x"54", -- $00a02
          x"55", -- $00a03
          x"52", -- $00a04
          x"4e", -- $00a05
          x"0a", -- $00a06
          x"0a", -- $00a07
          x"9f", -- $00a08
          x"9f", -- $00a09
          x"9d", -- $00a0a
          x"3c", -- $00a0b
          x"92", -- $00a0c
          x"3e", -- $00a0d
          x"92", -- $00a0e
          x"3f", -- $00a0f
          x"0a", -- $00a10
          x"20", -- $00a11
          x"4d", -- $00a12
          x"3d", -- $00a13
          x"91", -- $00a14
          x"53", -- $00a15
          x"48", -- $00a16
          x"49", -- $00a17
          x"46", -- $00a18
          x"54", -- $00a19
          x"91", -- $00a1a
          x"5a", -- $00a1b
          x"92", -- $00a1c
          x"58", -- $00a1d
          x"92", -- $00a1e
          x"43", -- $00a1f
          x"92", -- $00a20
          x"56", -- $00a21
          x"92", -- $00a22
          x"42", -- $00a23
          x"92", -- $00a24
          x"4e", -- $00a25
          x"92", -- $00a26
          x"4d", -- $00a27
          x"92", -- $00a28
          x"2c", -- $00a29
          x"92", -- $00a2a
          x"2e", -- $00a2b
          x"92", -- $00a2c
          x"2f", -- $00a2d
          x"92", -- $00a2e
          x"53", -- $00a2f
          x"48", -- $00a30
          x"49", -- $00a31
          x"46", -- $00a32
          x"54", -- $00a33
          x"91", -- $00a34
          x"55", -- $00a35
          x"50", -- $00a36
          x"0a", -- $00a37
          x"0a", -- $00a38
          x"9f", -- $00a39
          x"9f", -- $00a3a
          x"53", -- $00a3b
          x"50", -- $00a3c
          x"41", -- $00a3d
          x"43", -- $00a3e
          x"45", -- $00a3f
          x"0a", -- $00a40
          x"9f", -- $00a41
          x"9f", -- $00a42
          x"9f", -- $00a43
          x"9c", -- $00a44
          x"4c", -- $00a45
          x"45", -- $00a46
          x"46", -- $00a47
          x"54", -- $00a48
          x"20", -- $00a49
          x"44", -- $00a4a
          x"4f", -- $00a4b
          x"57", -- $00a4c
          x"4e", -- $00a4d
          x"20", -- $00a4e
          x"52", -- $00a4f
          x"47", -- $00a50
          x"48", -- $00a51
          x"54", -- $00a52
          x"0a", -- $00a53
          x"0a", -- $00a54
          x"0a", -- $00a55
          x"92", -- $00a56
          x"49", -- $00a57
          x"4e", -- $00a58
          x"46", -- $00a59
          x"4f", -- $00a5a
          x"52", -- $00a5b
          x"4d", -- $00a5c
          x"41", -- $00a5d
          x"54", -- $00a5e
          x"49", -- $00a5f
          x"4f", -- $00a60
          x"4e", -- $00a61
          x"41", -- $00a62
          x"4c", -- $00a63
          x"2d", -- $00a64
          x"54", -- $00a65
          x"45", -- $00a66
          x"58", -- $00a67
          x"54", -- $00a68
          x"2d", -- $00a69
          x"47", -- $00a6a
          x"4f", -- $00a6b
          x"45", -- $00a6c
          x"53", -- $00a6d
          x"2d", -- $00a6e
          x"48", -- $00a6f
          x"45", -- $00a70
          x"52", -- $00a71
          x"45", -- $00a72
          x"2e", -- $00a73
          x"2e", -- $00a74
          x"2e", -- $00a75
          x"2e", -- $00a76
          x"2e", -- $00a77
          x"2e", -- $00a78
          x"2e", -- $00a79
          x"0a", -- $00a7a
          x"92", -- $00a7b
          x"49", -- $00a7c
          x"4e", -- $00a7d
          x"46", -- $00a7e
          x"4f", -- $00a7f
          x"52", -- $00a80
          x"4d", -- $00a81
          x"41", -- $00a82
          x"54", -- $00a83
          x"49", -- $00a84
          x"4f", -- $00a85
          x"4e", -- $00a86
          x"41", -- $00a87
          x"4c", -- $00a88
          x"2d", -- $00a89
          x"54", -- $00a8a
          x"45", -- $00a8b
          x"58", -- $00a8c
          x"54", -- $00a8d
          x"2d", -- $00a8e
          x"47", -- $00a8f
          x"4f", -- $00a90
          x"45", -- $00a91
          x"53", -- $00a92
          x"2d", -- $00a93
          x"48", -- $00a94
          x"45", -- $00a95
          x"52", -- $00a96
          x"45", -- $00a97
          x"2e", -- $00a98
          x"2e", -- $00a99
          x"2e", -- $00a9a
          x"2e", -- $00a9b
          x"2e", -- $00a9c
          x"2e", -- $00a9d
          x"2e", -- $00a9e
          x"0a", -- $00a9f
          x"0a", -- $00aa0
          x"9f", -- $00aa1
          x"94", -- $00aa2
          x"fa", -- $00aa3
          x"f8", -- $00aa4
          x"0a", -- $00aa5
          x"93", -- $00aa6
          x"31", -- $00aa7
          x"92", -- $00aa8
          x"32", -- $00aa9
          x"92", -- $00aaa
          x"33", -- $00aab
          x"95", -- $00aac
          x"fb", -- $00aad
          x"f9", -- $00aae
          x"0a", -- $00aaf
          x"0a", -- $00ab0
          x"0a", -- $00ab1
          x"93", -- $00ab2
          x"34", -- $00ab3
          x"92", -- $00ab4
          x"35", -- $00ab5
          x"92", -- $00ab6
          x"36", -- $00ab7
          x"0a", -- $00ab8
          x"0a", -- $00ab9
          x"0a", -- $00aba
          x"93", -- $00abb
          x"37", -- $00abc
          x"92", -- $00abd
          x"38", -- $00abe
          x"92", -- $00abf
          x"39", -- $00ac0
          x"0a", -- $00ac1
          x"0a", -- $00ac2
          x"9f", -- $00ac3
          x"94", -- $00ac4
          x"fc", -- $00ac5
          x"fe", -- $00ac6
          x"0a", -- $00ac7
          x"93", -- $00ac8
          x"23", -- $00ac9
          x"92", -- $00aca
          x"30", -- $00acb
          x"92", -- $00acc
          x"2a", -- $00acd
          x"95", -- $00ace
          x"fd", -- $00acf
          x"ff", -- $00ad0
          x"0a", -- $00ad1
          x"0a", -- $00ad2
          x"0a", -- $00ad3
          x"00", -- $00ad4
          x"00", -- $00ad5
          x"00", -- $00ad6
          x"00", -- $00ad7
          x"00", -- $00ad8
          x"00", -- $00ad9
          x"00", -- $00ada
          x"00", -- $00adb
          x"00", -- $00adc
          x"00", -- $00add
          x"00", -- $00ade
          x"00", -- $00adf
          x"00", -- $00ae0
          x"00", -- $00ae1
          x"00", -- $00ae2
          x"00", -- $00ae3
          x"00", -- $00ae4
          x"00", -- $00ae5
          x"00", -- $00ae6
          x"00", -- $00ae7
          x"00", -- $00ae8
          x"00", -- $00ae9
          x"00", -- $00aea
          x"00", -- $00aeb
          x"00", -- $00aec
          x"00", -- $00aed
          x"00", -- $00aee
          x"00", -- $00aef
          x"00", -- $00af0
          x"00", -- $00af1
          x"00", -- $00af2
          x"00", -- $00af3
          x"00", -- $00af4
          x"00", -- $00af5
          x"00", -- $00af6
          x"00", -- $00af7
          x"00", -- $00af8
          x"00", -- $00af9
          x"00", -- $00afa
          x"00", -- $00afb
          x"00", -- $00afc
          x"00", -- $00afd
          x"00", -- $00afe
          x"00", -- $00aff
          x"00", -- $00b00
          x"00", -- $00b01
          x"00", -- $00b02
          x"00", -- $00b03
          x"00", -- $00b04
          x"00", -- $00b05
          x"00", -- $00b06
          x"00", -- $00b07
          x"00", -- $00b08
          x"00", -- $00b09
          x"00", -- $00b0a
          x"00", -- $00b0b
          x"00", -- $00b0c
          x"00", -- $00b0d
          x"00", -- $00b0e
          x"00", -- $00b0f
          x"00", -- $00b10
          x"00", -- $00b11
          x"00", -- $00b12
          x"00", -- $00b13
          x"00", -- $00b14
          x"00", -- $00b15
          x"00", -- $00b16
          x"00", -- $00b17
          x"00", -- $00b18
          x"00", -- $00b19
          x"00", -- $00b1a
          x"00", -- $00b1b
          x"00", -- $00b1c
          x"00", -- $00b1d
          x"00", -- $00b1e
          x"00", -- $00b1f
          x"00", -- $00b20
          x"00", -- $00b21
          x"00", -- $00b22
          x"00", -- $00b23
          x"00", -- $00b24
          x"00", -- $00b25
          x"00", -- $00b26
          x"00", -- $00b27
          x"00", -- $00b28
          x"00", -- $00b29
          x"00", -- $00b2a
          x"00", -- $00b2b
          x"00", -- $00b2c
          x"00", -- $00b2d
          x"00", -- $00b2e
          x"00", -- $00b2f
          x"00", -- $00b30
          x"00", -- $00b31
          x"00", -- $00b32
          x"00", -- $00b33
          x"00", -- $00b34
          x"00", -- $00b35
          x"00", -- $00b36
          x"00", -- $00b37
          x"00", -- $00b38
          x"00", -- $00b39
          x"00", -- $00b3a
          x"00", -- $00b3b
          x"00", -- $00b3c
          x"00", -- $00b3d
          x"00", -- $00b3e
          x"00", -- $00b3f
          x"00", -- $00b40
          x"00", -- $00b41
          x"00", -- $00b42
          x"00", -- $00b43
          x"00", -- $00b44
          x"00", -- $00b45
          x"00", -- $00b46
          x"00", -- $00b47
          x"00", -- $00b48
          x"00", -- $00b49
          x"00", -- $00b4a
          x"00", -- $00b4b
          x"00", -- $00b4c
          x"00", -- $00b4d
          x"00", -- $00b4e
          x"00", -- $00b4f
          x"00", -- $00b50
          x"00", -- $00b51
          x"00", -- $00b52
          x"00", -- $00b53
          x"00", -- $00b54
          x"00", -- $00b55
          x"00", -- $00b56
          x"00", -- $00b57
          x"00", -- $00b58
          x"00", -- $00b59
          x"00", -- $00b5a
          x"00", -- $00b5b
          x"00", -- $00b5c
          x"00", -- $00b5d
          x"00", -- $00b5e
          x"00", -- $00b5f
          x"00", -- $00b60
          x"00", -- $00b61
          x"00", -- $00b62
          x"00", -- $00b63
          x"00", -- $00b64
          x"00", -- $00b65
          x"00", -- $00b66
          x"00", -- $00b67
          x"00", -- $00b68
          x"00", -- $00b69
          x"00", -- $00b6a
          x"00", -- $00b6b
          x"00", -- $00b6c
          x"00", -- $00b6d
          x"00", -- $00b6e
          x"00", -- $00b6f
          x"00", -- $00b70
          x"00", -- $00b71
          x"00", -- $00b72
          x"00", -- $00b73
          x"00", -- $00b74
          x"00", -- $00b75
          x"00", -- $00b76
          x"00", -- $00b77
          x"00", -- $00b78
          x"00", -- $00b79
          x"00", -- $00b7a
          x"00", -- $00b7b
          x"00", -- $00b7c
          x"00", -- $00b7d
          x"00", -- $00b7e
          x"00", -- $00b7f
          x"00", -- $00b80
          x"00", -- $00b81
          x"00", -- $00b82
          x"00", -- $00b83
          x"00", -- $00b84
          x"00", -- $00b85
          x"00", -- $00b86
          x"00", -- $00b87
          x"00", -- $00b88
          x"00", -- $00b89
          x"00", -- $00b8a
          x"00", -- $00b8b
          x"00", -- $00b8c
          x"00", -- $00b8d
          x"00", -- $00b8e
          x"00", -- $00b8f
          x"00", -- $00b90
          x"00", -- $00b91
          x"00", -- $00b92
          x"00", -- $00b93
          x"00", -- $00b94
          x"00", -- $00b95
          x"00", -- $00b96
          x"00", -- $00b97
          x"00", -- $00b98
          x"00", -- $00b99
          x"00", -- $00b9a
          x"00", -- $00b9b
          x"00", -- $00b9c
          x"00", -- $00b9d
          x"00", -- $00b9e
          x"00", -- $00b9f
          x"00", -- $00ba0
          x"00", -- $00ba1
          x"00", -- $00ba2
          x"00", -- $00ba3
          x"00", -- $00ba4
          x"00", -- $00ba5
          x"00", -- $00ba6
          x"00", -- $00ba7
          x"00", -- $00ba8
          x"00", -- $00ba9
          x"00", -- $00baa
          x"00", -- $00bab
          x"00", -- $00bac
          x"00", -- $00bad
          x"00", -- $00bae
          x"00", -- $00baf
          x"00", -- $00bb0
          x"00", -- $00bb1
          x"00", -- $00bb2
          x"00", -- $00bb3
          x"00", -- $00bb4
          x"00", -- $00bb5
          x"00", -- $00bb6
          x"00", -- $00bb7
          x"00", -- $00bb8
          x"00", -- $00bb9
          x"00", -- $00bba
          x"00", -- $00bbb
          x"00", -- $00bbc
          x"00", -- $00bbd
          x"00", -- $00bbe
          x"00", -- $00bbf
          x"00", -- $00bc0
          x"00", -- $00bc1
          x"00", -- $00bc2
          x"00", -- $00bc3
          x"00", -- $00bc4
          x"00", -- $00bc5
          x"00", -- $00bc6
          x"00", -- $00bc7
          x"00", -- $00bc8
          x"00", -- $00bc9
          x"00", -- $00bca
          x"00", -- $00bcb
          x"00", -- $00bcc
          x"00", -- $00bcd
          x"00", -- $00bce
          x"00", -- $00bcf
          x"00", -- $00bd0
          x"00", -- $00bd1
          x"00", -- $00bd2
          x"00", -- $00bd3
          x"00", -- $00bd4
          x"00", -- $00bd5
          x"00", -- $00bd6
          x"00", -- $00bd7
          x"00", -- $00bd8
          x"00", -- $00bd9
          x"00", -- $00bda
          x"00", -- $00bdb
          x"00", -- $00bdc
          x"00", -- $00bdd
          x"00", -- $00bde
          x"00", -- $00bdf
          x"00", -- $00be0
          x"00", -- $00be1
          x"00", -- $00be2
          x"00", -- $00be3
          x"00", -- $00be4
          x"00", -- $00be5
          x"00", -- $00be6
          x"00", -- $00be7
          x"00", -- $00be8
          x"00", -- $00be9
          x"00", -- $00bea
          x"00", -- $00beb
          x"00", -- $00bec
          x"00", -- $00bed
          x"00", -- $00bee
          x"00", -- $00bef
          x"00", -- $00bf0
          x"00", -- $00bf1
          x"00", -- $00bf2
          x"00", -- $00bf3
          x"00", -- $00bf4
          x"00", -- $00bf5
          x"00", -- $00bf6
          x"00", -- $00bf7
          x"00", -- $00bf8
          x"00", -- $00bf9
          x"00", -- $00bfa
          x"00", -- $00bfb
          x"00", -- $00bfc
          x"00", -- $00bfd
          x"00", -- $00bfe
          x"00", -- $00bff
          x"00", -- $00c00
          x"00", -- $00c01
          x"00", -- $00c02
          x"00", -- $00c03
          x"00", -- $00c04
          x"00", -- $00c05
          x"00", -- $00c06
          x"00", -- $00c07
          x"00", -- $00c08
          x"00", -- $00c09
          x"00", -- $00c0a
          x"00", -- $00c0b
          x"00", -- $00c0c
          x"00", -- $00c0d
          x"00", -- $00c0e
          x"00", -- $00c0f
          x"00", -- $00c10
          x"00", -- $00c11
          x"00", -- $00c12
          x"00", -- $00c13
          x"00", -- $00c14
          x"00", -- $00c15
          x"00", -- $00c16
          x"00", -- $00c17
          x"00", -- $00c18
          x"00", -- $00c19
          x"00", -- $00c1a
          x"00", -- $00c1b
          x"00", -- $00c1c
          x"00", -- $00c1d
          x"00", -- $00c1e
          x"00", -- $00c1f
          x"00", -- $00c20
          x"00", -- $00c21
          x"00", -- $00c22
          x"00", -- $00c23
          x"00", -- $00c24
          x"00", -- $00c25
          x"00", -- $00c26
          x"00", -- $00c27
          x"00", -- $00c28
          x"00", -- $00c29
          x"00", -- $00c2a
          x"00", -- $00c2b
          x"00", -- $00c2c
          x"00", -- $00c2d
          x"00", -- $00c2e
          x"00", -- $00c2f
          x"00", -- $00c30
          x"00", -- $00c31
          x"00", -- $00c32
          x"00", -- $00c33
          x"00", -- $00c34
          x"00", -- $00c35
          x"00", -- $00c36
          x"00", -- $00c37
          x"00", -- $00c38
          x"00", -- $00c39
          x"00", -- $00c3a
          x"00", -- $00c3b
          x"00", -- $00c3c
          x"00", -- $00c3d
          x"00", -- $00c3e
          x"00", -- $00c3f
          x"00", -- $00c40
          x"00", -- $00c41
          x"00", -- $00c42
          x"00", -- $00c43
          x"00", -- $00c44
          x"00", -- $00c45
          x"00", -- $00c46
          x"00", -- $00c47
          x"00", -- $00c48
          x"00", -- $00c49
          x"00", -- $00c4a
          x"00", -- $00c4b
          x"00", -- $00c4c
          x"00", -- $00c4d
          x"00", -- $00c4e
          x"00", -- $00c4f
          x"00", -- $00c50
          x"00", -- $00c51
          x"00", -- $00c52
          x"00", -- $00c53
          x"00", -- $00c54
          x"00", -- $00c55
          x"00", -- $00c56
          x"00", -- $00c57
          x"00", -- $00c58
          x"00", -- $00c59
          x"00", -- $00c5a
          x"00", -- $00c5b
          x"00", -- $00c5c
          x"00", -- $00c5d
          x"00", -- $00c5e
          x"00", -- $00c5f
          x"00", -- $00c60
          x"00", -- $00c61
          x"00", -- $00c62
          x"00", -- $00c63
          x"00", -- $00c64
          x"00", -- $00c65
          x"00", -- $00c66
          x"00", -- $00c67
          x"00", -- $00c68
          x"00", -- $00c69
          x"00", -- $00c6a
          x"00", -- $00c6b
          x"00", -- $00c6c
          x"00", -- $00c6d
          x"00", -- $00c6e
          x"00", -- $00c6f
          x"00", -- $00c70
          x"00", -- $00c71
          x"00", -- $00c72
          x"00", -- $00c73
          x"00", -- $00c74
          x"00", -- $00c75
          x"00", -- $00c76
          x"00", -- $00c77
          x"00", -- $00c78
          x"00", -- $00c79
          x"00", -- $00c7a
          x"00", -- $00c7b
          x"00", -- $00c7c
          x"00", -- $00c7d
          x"00", -- $00c7e
          x"00", -- $00c7f
          x"00", -- $00c80
          x"00", -- $00c81
          x"00", -- $00c82
          x"00", -- $00c83
          x"00", -- $00c84
          x"00", -- $00c85
          x"00", -- $00c86
          x"00", -- $00c87
          x"00", -- $00c88
          x"00", -- $00c89
          x"00", -- $00c8a
          x"00", -- $00c8b
          x"00", -- $00c8c
          x"00", -- $00c8d
          x"00", -- $00c8e
          x"00", -- $00c8f
          x"00", -- $00c90
          x"00", -- $00c91
          x"00", -- $00c92
          x"00", -- $00c93
          x"00", -- $00c94
          x"00", -- $00c95
          x"00", -- $00c96
          x"00", -- $00c97
          x"00", -- $00c98
          x"00", -- $00c99
          x"00", -- $00c9a
          x"00", -- $00c9b
          x"00", -- $00c9c
          x"00", -- $00c9d
          x"00", -- $00c9e
          x"00", -- $00c9f
          x"00", -- $00ca0
          x"00", -- $00ca1
          x"00", -- $00ca2
          x"00", -- $00ca3
          x"00", -- $00ca4
          x"00", -- $00ca5
          x"00", -- $00ca6
          x"00", -- $00ca7
          x"00", -- $00ca8
          x"00", -- $00ca9
          x"00", -- $00caa
          x"00", -- $00cab
          x"00", -- $00cac
          x"00", -- $00cad
          x"00", -- $00cae
          x"00", -- $00caf
          x"00", -- $00cb0
          x"00", -- $00cb1
          x"00", -- $00cb2
          x"00", -- $00cb3
          x"00", -- $00cb4
          x"00", -- $00cb5
          x"00", -- $00cb6
          x"00", -- $00cb7
          x"00", -- $00cb8
          x"00", -- $00cb9
          x"00", -- $00cba
          x"00", -- $00cbb
          x"00", -- $00cbc
          x"00", -- $00cbd
          x"00", -- $00cbe
          x"00", -- $00cbf
          x"00", -- $00cc0
          x"00", -- $00cc1
          x"00", -- $00cc2
          x"00", -- $00cc3
          x"00", -- $00cc4
          x"00", -- $00cc5
          x"00", -- $00cc6
          x"00", -- $00cc7
          x"00", -- $00cc8
          x"00", -- $00cc9
          x"00", -- $00cca
          x"00", -- $00ccb
          x"00", -- $00ccc
          x"00", -- $00ccd
          x"00", -- $00cce
          x"00", -- $00ccf
          x"00", -- $00cd0
          x"00", -- $00cd1
          x"00", -- $00cd2
          x"00", -- $00cd3
          x"00", -- $00cd4
          x"00", -- $00cd5
          x"00", -- $00cd6
          x"00", -- $00cd7
          x"00", -- $00cd8
          x"00", -- $00cd9
          x"00", -- $00cda
          x"00", -- $00cdb
          x"00", -- $00cdc
          x"00", -- $00cdd
          x"00", -- $00cde
          x"00", -- $00cdf
          x"00", -- $00ce0
          x"00", -- $00ce1
          x"00", -- $00ce2
          x"00", -- $00ce3
          x"00", -- $00ce4
          x"00", -- $00ce5
          x"00", -- $00ce6
          x"00", -- $00ce7
          x"00", -- $00ce8
          x"00", -- $00ce9
          x"00", -- $00cea
          x"00", -- $00ceb
          x"00", -- $00cec
          x"00", -- $00ced
          x"00", -- $00cee
          x"00", -- $00cef
          x"00", -- $00cf0
          x"00", -- $00cf1
          x"00", -- $00cf2
          x"00", -- $00cf3
          x"00", -- $00cf4
          x"00", -- $00cf5
          x"00", -- $00cf6
          x"00", -- $00cf7
          x"00", -- $00cf8
          x"00", -- $00cf9
          x"00", -- $00cfa
          x"00", -- $00cfb
          x"00", -- $00cfc
          x"00", -- $00cfd
          x"00", -- $00cfe
          x"00", -- $00cff
          x"00", -- $00d00
          x"00", -- $00d01
          x"00", -- $00d02
          x"00", -- $00d03
          x"00", -- $00d04
          x"00", -- $00d05
          x"00", -- $00d06
          x"00", -- $00d07
          x"00", -- $00d08
          x"00", -- $00d09
          x"00", -- $00d0a
          x"00", -- $00d0b
          x"00", -- $00d0c
          x"00", -- $00d0d
          x"00", -- $00d0e
          x"00", -- $00d0f
          x"00", -- $00d10
          x"00", -- $00d11
          x"00", -- $00d12
          x"00", -- $00d13
          x"00", -- $00d14
          x"00", -- $00d15
          x"00", -- $00d16
          x"00", -- $00d17
          x"00", -- $00d18
          x"00", -- $00d19
          x"00", -- $00d1a
          x"00", -- $00d1b
          x"00", -- $00d1c
          x"00", -- $00d1d
          x"00", -- $00d1e
          x"00", -- $00d1f
          x"00", -- $00d20
          x"00", -- $00d21
          x"00", -- $00d22
          x"00", -- $00d23
          x"00", -- $00d24
          x"00", -- $00d25
          x"00", -- $00d26
          x"00", -- $00d27
          x"00", -- $00d28
          x"00", -- $00d29
          x"00", -- $00d2a
          x"00", -- $00d2b
          x"00", -- $00d2c
          x"00", -- $00d2d
          x"00", -- $00d2e
          x"00", -- $00d2f
          x"00", -- $00d30
          x"00", -- $00d31
          x"00", -- $00d32
          x"00", -- $00d33
          x"00", -- $00d34
          x"00", -- $00d35
          x"00", -- $00d36
          x"00", -- $00d37
          x"00", -- $00d38
          x"00", -- $00d39
          x"00", -- $00d3a
          x"00", -- $00d3b
          x"00", -- $00d3c
          x"00", -- $00d3d
          x"00", -- $00d3e
          x"00", -- $00d3f
          x"00", -- $00d40
          x"00", -- $00d41
          x"00", -- $00d42
          x"00", -- $00d43
          x"00", -- $00d44
          x"00", -- $00d45
          x"00", -- $00d46
          x"00", -- $00d47
          x"00", -- $00d48
          x"00", -- $00d49
          x"00", -- $00d4a
          x"00", -- $00d4b
          x"00", -- $00d4c
          x"00", -- $00d4d
          x"00", -- $00d4e
          x"00", -- $00d4f
          x"00", -- $00d50
          x"00", -- $00d51
          x"00", -- $00d52
          x"00", -- $00d53
          x"00", -- $00d54
          x"00", -- $00d55
          x"00", -- $00d56
          x"00", -- $00d57
          x"00", -- $00d58
          x"00", -- $00d59
          x"00", -- $00d5a
          x"00", -- $00d5b
          x"00", -- $00d5c
          x"00", -- $00d5d
          x"00", -- $00d5e
          x"00", -- $00d5f
          x"00", -- $00d60
          x"00", -- $00d61
          x"00", -- $00d62
          x"00", -- $00d63
          x"00", -- $00d64
          x"00", -- $00d65
          x"00", -- $00d66
          x"00", -- $00d67
          x"00", -- $00d68
          x"00", -- $00d69
          x"00", -- $00d6a
          x"00", -- $00d6b
          x"00", -- $00d6c
          x"00", -- $00d6d
          x"00", -- $00d6e
          x"00", -- $00d6f
          x"00", -- $00d70
          x"00", -- $00d71
          x"00", -- $00d72
          x"00", -- $00d73
          x"00", -- $00d74
          x"00", -- $00d75
          x"00", -- $00d76
          x"00", -- $00d77
          x"00", -- $00d78
          x"00", -- $00d79
          x"00", -- $00d7a
          x"00", -- $00d7b
          x"00", -- $00d7c
          x"00", -- $00d7d
          x"00", -- $00d7e
          x"00", -- $00d7f
          x"00", -- $00d80
          x"00", -- $00d81
          x"00", -- $00d82
          x"00", -- $00d83
          x"00", -- $00d84
          x"00", -- $00d85
          x"00", -- $00d86
          x"00", -- $00d87
          x"00", -- $00d88
          x"00", -- $00d89
          x"00", -- $00d8a
          x"00", -- $00d8b
          x"00", -- $00d8c
          x"00", -- $00d8d
          x"00", -- $00d8e
          x"00", -- $00d8f
          x"00", -- $00d90
          x"00", -- $00d91
          x"00", -- $00d92
          x"00", -- $00d93
          x"00", -- $00d94
          x"00", -- $00d95
          x"00", -- $00d96
          x"00", -- $00d97
          x"00", -- $00d98
          x"00", -- $00d99
          x"00", -- $00d9a
          x"00", -- $00d9b
          x"00", -- $00d9c
          x"00", -- $00d9d
          x"00", -- $00d9e
          x"00", -- $00d9f
          x"00", -- $00da0
          x"00", -- $00da1
          x"00", -- $00da2
          x"00", -- $00da3
          x"00", -- $00da4
          x"00", -- $00da5
          x"00", -- $00da6
          x"00", -- $00da7
          x"00", -- $00da8
          x"00", -- $00da9
          x"00", -- $00daa
          x"00", -- $00dab
          x"00", -- $00dac
          x"00", -- $00dad
          x"00", -- $00dae
          x"00", -- $00daf
          x"00", -- $00db0
          x"00", -- $00db1
          x"00", -- $00db2
          x"00", -- $00db3
          x"00", -- $00db4
          x"00", -- $00db5
          x"00", -- $00db6
          x"00", -- $00db7
          x"00", -- $00db8
          x"00", -- $00db9
          x"00", -- $00dba
          x"00", -- $00dbb
          x"00", -- $00dbc
          x"00", -- $00dbd
          x"00", -- $00dbe
          x"00", -- $00dbf
          x"00", -- $00dc0
          x"00", -- $00dc1
          x"00", -- $00dc2
          x"00", -- $00dc3
          x"00", -- $00dc4
          x"00", -- $00dc5
          x"00", -- $00dc6
          x"00", -- $00dc7
          x"00", -- $00dc8
          x"00", -- $00dc9
          x"00", -- $00dca
          x"00", -- $00dcb
          x"00", -- $00dcc
          x"00", -- $00dcd
          x"00", -- $00dce
          x"00", -- $00dcf
          x"00", -- $00dd0
          x"00", -- $00dd1
          x"00", -- $00dd2
          x"00", -- $00dd3
          x"00", -- $00dd4
          x"00", -- $00dd5
          x"00", -- $00dd6
          x"00", -- $00dd7
          x"00", -- $00dd8
          x"00", -- $00dd9
          x"00", -- $00dda
          x"00", -- $00ddb
          x"00", -- $00ddc
          x"00", -- $00ddd
          x"00", -- $00dde
          x"00", -- $00ddf
          x"00", -- $00de0
          x"00", -- $00de1
          x"00", -- $00de2
          x"00", -- $00de3
          x"00", -- $00de4
          x"00", -- $00de5
          x"00", -- $00de6
          x"00", -- $00de7
          x"00", -- $00de8
          x"00", -- $00de9
          x"00", -- $00dea
          x"00", -- $00deb
          x"00", -- $00dec
          x"00", -- $00ded
          x"00", -- $00dee
          x"00", -- $00def
          x"00", -- $00df0
          x"00", -- $00df1
          x"00", -- $00df2
          x"00", -- $00df3
          x"00", -- $00df4
          x"00", -- $00df5
          x"00", -- $00df6
          x"00", -- $00df7
          x"00", -- $00df8
          x"00", -- $00df9
          x"00", -- $00dfa
          x"00", -- $00dfb
          x"00", -- $00dfc
          x"00", -- $00dfd
          x"00", -- $00dfe
          x"00", -- $00dff
          x"7e", -- $00e00
          x"02", -- $00e01
          x"7e", -- $00e02
          x"04", -- $00e03
          x"08", -- $00e04
          x"30", -- $00e05
          x"00", -- $00e06
          x"00", -- $00e07
          x"00", -- $00e08
          x"00", -- $00e09
          x"7c", -- $00e0a
          x"1e", -- $00e0b
          x"10", -- $00e0c
          x"10", -- $00e0d
          x"20", -- $00e0e
          x"00", -- $00e0f
          x"00", -- $00e10
          x"04", -- $00e11
          x"0c", -- $00e12
          x"18", -- $00e13
          x"68", -- $00e14
          x"08", -- $00e15
          x"08", -- $00e16
          x"00", -- $00e17
          x"00", -- $00e18
          x"10", -- $00e19
          x"7c", -- $00e1a
          x"44", -- $00e1b
          x"44", -- $00e1c
          x"08", -- $00e1d
          x"10", -- $00e1e
          x"00", -- $00e1f
          x"00", -- $00e20
          x"00", -- $00e21
          x"7c", -- $00e22
          x"10", -- $00e23
          x"10", -- $00e24
          x"7c", -- $00e25
          x"00", -- $00e26
          x"00", -- $00e27
          x"00", -- $00e28
          x"08", -- $00e29
          x"7e", -- $00e2a
          x"18", -- $00e2b
          x"18", -- $00e2c
          x"68", -- $00e2d
          x"18", -- $00e2e
          x"00", -- $00e2f
          x"00", -- $00e30
          x"20", -- $00e31
          x"1e", -- $00e32
          x"74", -- $00e33
          x"14", -- $00e34
          x"08", -- $00e35
          x"08", -- $00e36
          x"00", -- $00e37
          x"00", -- $00e38
          x"00", -- $00e39
          x"78", -- $00e3a
          x"08", -- $00e3b
          x"08", -- $00e3c
          x"7e", -- $00e3d
          x"00", -- $00e3e
          x"00", -- $00e3f
          x"7e", -- $00e40
          x"04", -- $00e41
          x"34", -- $00e42
          x"0c", -- $00e43
          x"36", -- $00e44
          x"44", -- $00e45
          x"00", -- $00e46
          x"00", -- $00e47
          x"00", -- $00e48
          x"00", -- $00e49
          x"74", -- $00e4a
          x"54", -- $00e4b
          x"2c", -- $00e4c
          x"08", -- $00e4d
          x"30", -- $00e4e
          x"00", -- $00e4f
          x"40", -- $00e50
          x"22", -- $00e51
          x"02", -- $00e52
          x"06", -- $00e53
          x"08", -- $00e54
          x"70", -- $00e55
          x"00", -- $00e56
          x"00", -- $00e57
          x"7f", -- $00e58
          x"02", -- $00e59
          x"0c", -- $00e5a
          x"08", -- $00e5b
          x"08", -- $00e5c
          x"10", -- $00e5d
          x"30", -- $00e5e
          x"00", -- $00e5f
          x"06", -- $00e60
          x"04", -- $00e61
          x"08", -- $00e62
          x"38", -- $00e63
          x"48", -- $00e64
          x"08", -- $00e65
          x"08", -- $00e66
          x"00", -- $00e67
          x"10", -- $00e68
          x"7e", -- $00e69
          x"42", -- $00e6a
          x"42", -- $00e6b
          x"04", -- $00e6c
          x"0c", -- $00e6d
          x"18", -- $00e6e
          x"00", -- $00e6f
          x"00", -- $00e70
          x"3e", -- $00e71
          x"08", -- $00e72
          x"08", -- $00e73
          x"08", -- $00e74
          x"7f", -- $00e75
          x"00", -- $00e76
          x"00", -- $00e77
          x"04", -- $00e78
          x"3f", -- $00e79
          x"0c", -- $00e7a
          x"0c", -- $00e7b
          x"14", -- $00e7c
          x"24", -- $00e7d
          x"4c", -- $00e7e
          x"00", -- $00e7f
          x"10", -- $00e80
          x"7e", -- $00e81
          x"12", -- $00e82
          x"12", -- $00e83
          x"22", -- $00e84
          x"4e", -- $00e85
          x"00", -- $00e86
          x"00", -- $00e87
          x"10", -- $00e88
          x"0e", -- $00e89
          x"78", -- $00e8a
          x"0b", -- $00e8b
          x"7c", -- $00e8c
          x"0c", -- $00e8d
          x"04", -- $00e8e
          x"00", -- $00e8f
          x"18", -- $00e90
          x"1e", -- $00e91
          x"32", -- $00e92
          x"62", -- $00e93
          x"04", -- $00e94
          x"08", -- $00e95
          x"30", -- $00e96
          x"00", -- $00e97
          x"10", -- $00e98
          x"3f", -- $00e99
          x"64", -- $00e9a
          x"44", -- $00e9b
          x"08", -- $00e9c
          x"08", -- $00e9d
          x"10", -- $00e9e
          x"00", -- $00e9f
          x"00", -- $00ea0
          x"7c", -- $00ea1
          x"04", -- $00ea2
          x"04", -- $00ea3
          x"04", -- $00ea4
          x"7c", -- $00ea5
          x"00", -- $00ea6
          x"00", -- $00ea7
          x"22", -- $00ea8
          x"22", -- $00ea9
          x"7f", -- $00eaa
          x"22", -- $00eab
          x"22", -- $00eac
          x"04", -- $00ead
          x"08", -- $00eae
          x"00", -- $00eaf
          x"20", -- $00eb0
          x"10", -- $00eb1
          x"63", -- $00eb2
          x"06", -- $00eb3
          x"0c", -- $00eb4
          x"30", -- $00eb5
          x"00", -- $00eb6
          x"00", -- $00eb7
          x"3e", -- $00eb8
          x"04", -- $00eb9
          x"08", -- $00eba
          x"1c", -- $00ebb
          x"32", -- $00ebc
          x"43", -- $00ebd
          x"00", -- $00ebe
          x"00", -- $00ebf
          x"10", -- $00ec0
          x"12", -- $00ec1
          x"7f", -- $00ec2
          x"14", -- $00ec3
          x"10", -- $00ec4
          x"1e", -- $00ec5
          x"00", -- $00ec6
          x"00", -- $00ec7
          x"42", -- $00ec8
          x"62", -- $00ec9
          x"22", -- $00eca
          x"04", -- $00ecb
          x"0c", -- $00ecc
          x"08", -- $00ecd
          x"30", -- $00ece
          x"00", -- $00ecf
          x"10", -- $00ed0
          x"3c", -- $00ed1
          x"26", -- $00ed2
          x"54", -- $00ed3
          x"0c", -- $00ed4
          x"18", -- $00ed5
          x"20", -- $00ed6
          x"00", -- $00ed7
          x"1e", -- $00ed8
          x"28", -- $00ed9
          x"7f", -- $00eda
          x"08", -- $00edb
          x"08", -- $00edc
          x"10", -- $00edd
          x"30", -- $00ede
          x"00", -- $00edf
          x"3e", -- $00ee0
          x"00", -- $00ee1
          x"7f", -- $00ee2
          x"08", -- $00ee3
          x"08", -- $00ee4
          x"08", -- $00ee5
          x"10", -- $00ee6
          x"00", -- $00ee7
          x"08", -- $00ee8
          x"1c", -- $00ee9
          x"26", -- $00eea
          x"0c", -- $00eeb
          x"3b", -- $00eec
          x"48", -- $00eed
          x"08", -- $00eee
          x"00", -- $00eef
          x"08", -- $00ef0
          x"08", -- $00ef1
          x"7f", -- $00ef2
          x"08", -- $00ef3
          x"08", -- $00ef4
          x"18", -- $00ef5
          x"30", -- $00ef6
          x"00", -- $00ef7
          x"08", -- $00ef8
          x"7f", -- $00ef9
          x"08", -- $00efa
          x"2a", -- $00efb
          x"2b", -- $00efc
          x"49", -- $00efd
          x"08", -- $00efe
          x"00", -- $00eff
          x"00", -- $00f00
          x"00", -- $00f01
          x"00", -- $00f02
          x"00", -- $00f03
          x"00", -- $00f04
          x"00", -- $00f05
          x"00", -- $00f06
          x"00", -- $00f07
          x"00", -- $00f08
          x"00", -- $00f09
          x"00", -- $00f0a
          x"00", -- $00f0b
          x"00", -- $00f0c
          x"00", -- $00f0d
          x"00", -- $00f0e
          x"00", -- $00f0f
          x"00", -- $00f10
          x"00", -- $00f11
          x"00", -- $00f12
          x"00", -- $00f13
          x"00", -- $00f14
          x"00", -- $00f15
          x"00", -- $00f16
          x"00", -- $00f17
          x"00", -- $00f18
          x"00", -- $00f19
          x"00", -- $00f1a
          x"00", -- $00f1b
          x"00", -- $00f1c
          x"00", -- $00f1d
          x"00", -- $00f1e
          x"00", -- $00f1f
          x"00", -- $00f20
          x"00", -- $00f21
          x"00", -- $00f22
          x"00", -- $00f23
          x"00", -- $00f24
          x"00", -- $00f25
          x"00", -- $00f26
          x"00", -- $00f27
          x"00", -- $00f28
          x"00", -- $00f29
          x"00", -- $00f2a
          x"00", -- $00f2b
          x"00", -- $00f2c
          x"00", -- $00f2d
          x"00", -- $00f2e
          x"00", -- $00f2f
          x"00", -- $00f30
          x"00", -- $00f31
          x"00", -- $00f32
          x"00", -- $00f33
          x"00", -- $00f34
          x"00", -- $00f35
          x"00", -- $00f36
          x"00", -- $00f37
          x"00", -- $00f38
          x"00", -- $00f39
          x"00", -- $00f3a
          x"00", -- $00f3b
          x"00", -- $00f3c
          x"00", -- $00f3d
          x"00", -- $00f3e
          x"00", -- $00f3f
          x"00", -- $00f40
          x"00", -- $00f41
          x"00", -- $00f42
          x"00", -- $00f43
          x"00", -- $00f44
          x"00", -- $00f45
          x"00", -- $00f46
          x"00", -- $00f47
          x"00", -- $00f48
          x"00", -- $00f49
          x"00", -- $00f4a
          x"00", -- $00f4b
          x"00", -- $00f4c
          x"00", -- $00f4d
          x"00", -- $00f4e
          x"00", -- $00f4f
          x"00", -- $00f50
          x"00", -- $00f51
          x"00", -- $00f52
          x"00", -- $00f53
          x"00", -- $00f54
          x"00", -- $00f55
          x"00", -- $00f56
          x"00", -- $00f57
          x"00", -- $00f58
          x"00", -- $00f59
          x"00", -- $00f5a
          x"00", -- $00f5b
          x"00", -- $00f5c
          x"00", -- $00f5d
          x"00", -- $00f5e
          x"00", -- $00f5f
          x"00", -- $00f60
          x"00", -- $00f61
          x"00", -- $00f62
          x"00", -- $00f63
          x"00", -- $00f64
          x"00", -- $00f65
          x"00", -- $00f66
          x"00", -- $00f67
          x"00", -- $00f68
          x"00", -- $00f69
          x"00", -- $00f6a
          x"00", -- $00f6b
          x"00", -- $00f6c
          x"00", -- $00f6d
          x"00", -- $00f6e
          x"00", -- $00f6f
          x"00", -- $00f70
          x"00", -- $00f71
          x"00", -- $00f72
          x"00", -- $00f73
          x"00", -- $00f74
          x"00", -- $00f75
          x"00", -- $00f76
          x"00", -- $00f77
          x"00", -- $00f78
          x"00", -- $00f79
          x"00", -- $00f7a
          x"00", -- $00f7b
          x"00", -- $00f7c
          x"00", -- $00f7d
          x"00", -- $00f7e
          x"00", -- $00f7f
          x"00", -- $00f80
          x"00", -- $00f81
          x"00", -- $00f82
          x"00", -- $00f83
          x"00", -- $00f84
          x"00", -- $00f85
          x"00", -- $00f86
          x"00", -- $00f87
          x"00", -- $00f88
          x"00", -- $00f89
          x"00", -- $00f8a
          x"00", -- $00f8b
          x"00", -- $00f8c
          x"00", -- $00f8d
          x"00", -- $00f8e
          x"00", -- $00f8f
          x"00", -- $00f90
          x"00", -- $00f91
          x"00", -- $00f92
          x"00", -- $00f93
          x"00", -- $00f94
          x"00", -- $00f95
          x"00", -- $00f96
          x"00", -- $00f97
          x"00", -- $00f98
          x"00", -- $00f99
          x"00", -- $00f9a
          x"00", -- $00f9b
          x"00", -- $00f9c
          x"00", -- $00f9d
          x"00", -- $00f9e
          x"00", -- $00f9f
          x"00", -- $00fa0
          x"00", -- $00fa1
          x"00", -- $00fa2
          x"00", -- $00fa3
          x"00", -- $00fa4
          x"00", -- $00fa5
          x"00", -- $00fa6
          x"00", -- $00fa7
          x"00", -- $00fa8
          x"00", -- $00fa9
          x"00", -- $00faa
          x"00", -- $00fab
          x"00", -- $00fac
          x"00", -- $00fad
          x"00", -- $00fae
          x"00", -- $00faf
          x"00", -- $00fb0
          x"00", -- $00fb1
          x"00", -- $00fb2
          x"00", -- $00fb3
          x"00", -- $00fb4
          x"00", -- $00fb5
          x"00", -- $00fb6
          x"00", -- $00fb7
          x"00", -- $00fb8
          x"00", -- $00fb9
          x"00", -- $00fba
          x"00", -- $00fbb
          x"00", -- $00fbc
          x"00", -- $00fbd
          x"00", -- $00fbe
          x"00", -- $00fbf
          x"00", -- $00fc0
          x"00", -- $00fc1
          x"00", -- $00fc2
          x"00", -- $00fc3
          x"00", -- $00fc4
          x"00", -- $00fc5
          x"00", -- $00fc6
          x"00", -- $00fc7
          x"00", -- $00fc8
          x"00", -- $00fc9
          x"00", -- $00fca
          x"00", -- $00fcb
          x"00", -- $00fcc
          x"00", -- $00fcd
          x"00", -- $00fce
          x"00", -- $00fcf
          x"00", -- $00fd0
          x"00", -- $00fd1
          x"00", -- $00fd2
          x"00", -- $00fd3
          x"00", -- $00fd4
          x"00", -- $00fd5
          x"00", -- $00fd6
          x"00", -- $00fd7
          x"00", -- $00fd8
          x"00", -- $00fd9
          x"00", -- $00fda
          x"00", -- $00fdb
          x"00", -- $00fdc
          x"00", -- $00fdd
          x"00", -- $00fde
          x"00", -- $00fdf
          x"00", -- $00fe0
          x"00", -- $00fe1
          x"00", -- $00fe2
          x"00", -- $00fe3
          x"00", -- $00fe4
          x"00", -- $00fe5
          x"00", -- $00fe6
          x"00", -- $00fe7
          x"00", -- $00fe8
          x"00", -- $00fe9
          x"00", -- $00fea
          x"00", -- $00feb
          x"00", -- $00fec
          x"00", -- $00fed
          x"00", -- $00fee
          x"00", -- $00fef
          x"00", -- $00ff0
          x"00", -- $00ff1
          x"00", -- $00ff2
          x"00", -- $00ff3
          x"00", -- $00ff4
          x"00", -- $00ff5
          x"00", -- $00ff6
          x"00", -- $00ff7
          x"00", -- $00ff8
          x"00", -- $00ff9
          x"00", -- $00ffa
          x"00", -- $00ffb
          x"00", -- $00ffc
          x"55", -- $00ffd
          x"0a", -- $00ffe
          x"0f"); -- $00fff
  shared variable ram : ram_t := initram;
begin

--process for read and write operation.
  PROCESS(Clk,write_count,no_write_count)
  BEGIN
    writes <= write_count;
    no_writes <= no_write_count;
    data_o <= ram(address);
    if(rising_edge(Clk)) then 
      if we /= '0' then
        write_count <= write_count + 1;        
        ram(address) := data_i;
      else
        no_write_count <= no_write_count + 1;        
      end if;
    end if;
  END PROCESS;

end Behavioral;
